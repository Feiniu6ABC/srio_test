

//protect begin

//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/common/srio_gen2_v4_1_16_cfg_axi.v#3 $
//----------------------------------------------------------------------
//
// CFG_AXI
// Description:
// This module contains the configuration register interface used for
// each core.
//
// It uses an AXI-Lite interface to the Configuration Fabric, and has a
// core interface for transfer of control and status information.
//
// No clock relationship between the cfg_clk and the core's clock is
// assumed.
//
// Hierarchy:
// LOG_TOP
//    |______LOG_CFG_TOP
//              |______CFG_AXI <-- this module
//              |______LOG_CFG_REG
// BUF_TOP
//    |______BUF_CFG_TOP
//              |______CFG_AXI <-- this module
//              |______BUF_CFG_REG
// PHY_TOP
//    |______PHY_CFG_TOP
//              |______CFG_AXI <-- this module
//              |______PHY_CFG_REG
// ---------------------------------------------------------------------
`timescale 1ps/1ps

// ------------------------------------------------
// below attribute is added to supress the synthesis warnings in vivado tool 8:3332
(* DowngradeIPIdentifiedWarnings="yes" *)
// ------------------------------------------------

module srio_gen2_v4_1_16_cfg_axi
  #(
    parameter TCQ   = 100)
  (
    // {{{ Port Declarations ---------------
    // System Signals
    input             core_clk,           // Core interface clock (phy_clk for PHY, etc.)
    input             cfg_clk,            // CFG Interface user clock
    input             cfg_rst,            // Reset for CFG clk domain

    // Configuration Fabric Interface
    input             CF_awvalid,         // Write Address Valid
    output reg        CCA_awready,        // Write Address Port Ready
    input      [23:0] CF_awaddr,          // Write Address
    input             CF_wvalid,          // Write Data Valid
    output reg        CCA_wready,         // Write Data Port Ready
    input      [31:0] CF_wdata,           // Write Data
    input      [ 3:0] CF_wstrb,           // Write Data Byte Enables
    output reg        CCA_bvalid,         // Write Response Valid
    input             CF_bready,          // Write Response Fabric Ready
    input             CF_arvalid,         // Read Address Valid
    output reg        CCA_arready,        // Read Address Port Ready
    input      [23:0] CF_araddr,          // Read Address
    output reg        CCA_rvalid,         // Read Response Valid
    input             CF_rready,          // Read Response Fabric Ready
    output reg [31:0] CCA_rdata,          // Read Data

    // Configuration Register Interface
    output reg        CCA_sync_cfg_rst,   // cfg_rst sync'ed to core_clk
    output reg [23:0] CCA_cfg_waddr,      // Write Address
    output reg [31:0] CCA_cfg_wdata,      // Write Data
    output reg [3:0]  CCA_cfg_wstrb,      // Write Data Byte Enables
    output reg        CCA_sync_we,        // Synchronized write enable
    output reg [23:0] CCA_cfg_raddr,      // Read Address
    output reg        CCA_sync_re,        // Synchronized Read Enable
    input      [31:0] CC_core_rdata       // Read Data
    // }}} End Port Declarations -----------
  );
  // {{{ Wire Declarations -----------------
  reg           cfg_rst_q;                // registered version of cfg_rst (cfg_clk domain)
  reg           cfg_rst_qq;               // registered version of cfg_rst_q to set readys to 1
  reg [1:0]     cfg_rst_sync;             // synchronization reg for cfg_rst in core_clk domain
  reg [1:0]     cfg_rst_resync;           // synchronization reg for CCA_sync_cfg_rst back to cfg_clk domain
  reg           cfg_rst_resync_q;         // registered version of cfg_rst_resync[1] used to detect falling edge
  reg           set_ready_post_reset;     // Set readys after reset is synchronized back to core_clk
  wire          wdata_active;             // write data xfer in progress (wvalid AND wready)
  reg           got_wdata;                // write data and strobe captured from Config Fabric
  wire          waddr_active;             // write address xfer in progress (awvalid AND awready)
  reg           got_waddr;                // write address captured from Config Fabric
  wire          set_we;                   // write info received (got_wdata AND got_waddr)
  wire          raddr_active;             // read address xfer in progress (arvalid AND arready)
  wire          rresp_active;             // read response xfer in progress (rvalid AND rready)
  reg           wsync_cfg_req = 0;        // cfg_clk domain register stage for write synchronization
  (* shreg_extract = "no" *)              // prevent the tools from inferring a shift register on synchronizer
  reg           wsync_core_q = 0;         // core_clk domain register stage for write synchronization
  (* shreg_extract = "no" *)
  reg           bsync_core_req = 0;       // core_clk domain register stage for write synchronization
  (* shreg_extract = "no" *)
  reg           bsync_cfg_q = 0;          // cfg_clk domain register stage for write synchronization
  (* shreg_extract = "no" *)
  reg           bsync_cfg_done = 0;       // write is complete and it is safe to accept new data/address
  reg           bsync_cfg_hold_done = 0;  // hold the above signal until write response accepted by config fabric
  wire          bsync_cfg_complete;       // OR of the two previous signals, used to release readys
  reg           arsync_cfg_req = 0;       // cfg_clk domain register stage for read address synchronization
  (* shreg_extract = "no" *)
  reg           arsync_core_q = 0;        // core_clk domain register stage for read address synchronization
  (* shreg_extract = "no" *)
  reg           rsync_core_req = 0;       // start sync back to know when read data can be sampled for resp
  (* shreg_extract = "no" *)
  reg           rsync_cfg_q = 0;          // cfg_clk domain register stage for read response synchronization
  (* shreg_extract = "no" *)
  reg           rsync_cfg_done = 0;       // read response synchronization done - safe to sample read data
  // }}} End Wire Declarations -------------

  // {{{ Reset Fanout Control --------------
  // Register cfg_rst before use (set asynchronously for immediate
  // availability)
  always @(posedge cfg_clk or posedge cfg_rst) begin
    if (cfg_rst) begin
      cfg_rst_q       <=  #TCQ 1'b1;
    end else begin
      cfg_rst_q       <=  #TCQ 1'b0;
    end
  end

  // Register reset again so that readys can be set back to 1.
  always @(posedge cfg_clk) begin
    cfg_rst_qq        <=  #TCQ cfg_rst_q;
  end

  // Synchronize cfg_aresetn to core_clk domain.
  // Will assert for multiple core_clk cycles and deassert synchronously.
  always @(posedge core_clk or posedge cfg_rst) begin
    if (cfg_rst) begin
      cfg_rst_sync        <=  #TCQ 2'b11;
      CCA_sync_cfg_rst    <=  #TCQ 1'b1;
    end else begin
      cfg_rst_sync        <=  #TCQ {cfg_rst_sync[0], 1'b0};
      CCA_sync_cfg_rst    <=  #TCQ  cfg_rst_sync[1];
    end
  end
  

  // Synchronize reset back to cfg_clk domain
  always @(posedge cfg_clk or posedge CCA_sync_cfg_rst) begin
    if (CCA_sync_cfg_rst) begin
      cfg_rst_resync        <= #TCQ 2'b11;
    end else begin
      cfg_rst_resync        <= #TCQ {cfg_rst_resync[0], 1'b0};
    end
  end
  always @(posedge cfg_clk) begin
    cfg_rst_resync_q      <= #TCQ cfg_rst_resync[1];
    set_ready_post_reset  <= #TCQ cfg_rst_resync_q && !cfg_rst_resync[1];
  end

  // }}} End Reset Fanout Control ----------

  // {{{ Wait for Write Data/Address -------
  // This block controls the Write Address and Write Data channels on the
  // AXI-Lite interface to the Configuration Fabric.
  // It must hold off the write until both address and data have been received.

  //*COVERPOINT*
  //(cp_simultaneous_waddr_and_wdata): Received Write Address and Data at the same time
  //(cp_wdata_before_waddr): Received Write Data before Address
  //(cp_waddr_before_wdata): Received Write Address before Data

  // Create signals to indicate transfer of data/address in progress
  assign wdata_active = CF_wvalid  && CCA_wready;
  assign waddr_active = CF_awvalid && CCA_awready;

  //*ASSERTION*
  //(ap_set_we_asserted_with_waddr_active): waddr_active should not assert while set_we is high

  // Indicate that write address was received
  always @(posedge cfg_clk) begin
    if (cfg_rst_q) begin
      got_waddr       <= #TCQ 1'b0;
    end else if (waddr_active) begin
      got_waddr       <= #TCQ 1'b1;
    end else if (set_we) begin
      got_waddr       <= #TCQ 1'b0;
    end
  end

  //*ASSERTION*
  //(ap_set_we_asserted_with_wdata_active): wdata_active should not assert while set_we is high

  // Indicate that write data (and strobe) received
  always @(posedge cfg_clk) begin
    if (cfg_rst_q) begin
      got_wdata       <= #TCQ 1'b0;
    end else if (wdata_active) begin
      got_wdata       <= #TCQ 1'b1;
    end else if (set_we) begin
      got_wdata       <= #TCQ 1'b0;
    end
  end

  // Create signal to start write sync process once both write data and address
  // are available.
  // Can remove a cycle of latency by looking at w<data/addr>_active signals, but that uses unreg inputs
  //*ASSERTION*
  //(ap_waddr_wdata_cnt_mismatch): Should accept equal number of waddrs and wdatas
  //*COVERPOINT*
  //(cp_reset_set_we): Reset on same cycle as set_we asserts
  assign set_we = (got_waddr && got_wdata);

  // Capture write address from Config Fabric
  // No reset needed for waddr_q - it's a don't care until a valid address is
  // received.
  //*ASSERTION*
  //(ap_waddr_sampled_incorrectly): cfg_waddr should be the same as the accepted address when sync_we asserts
  always @(posedge cfg_clk) begin
    if (CCA_awready) begin
      CCA_cfg_waddr   <= #TCQ {CF_awaddr[23:2], 2'b0}; // Tying off lower bits results in less address decode logic
    end
  end

  // Capture write data and strobe from Config Fabric
  // No reset needed for wdata_q or wstrb_q - they're don't cares until valid
  // information is received.
  //*ASSERTION*
  //(ap_wdata_sampled_incorrectly): cfg_wdata should be the same as the accepted data when sync_we asserts
  //(ap_wstrb_sampled_incorrectly): cfg_wstrb should be the same as the accepted strobe when sync_we asserts
  always @(posedge cfg_clk) begin
    if (CCA_wready) begin
      CCA_cfg_wdata   <= #TCQ CF_wdata;
      CCA_cfg_wstrb   <= #TCQ CF_wstrb;
    end
  end

  // Create awready output - hold low after addr is captured until write completes
  // IP Checklist violation - Using unreg inputs (awvalid as part of waddr_active)
  always @(posedge cfg_clk) begin
    if (cfg_rst_q) begin
      CCA_awready     <= #TCQ 1'b0;
    end else if (set_ready_post_reset) begin              // Set to 1 after reset
      CCA_awready     <= #TCQ 1'b1;
    end else if (waddr_active || got_waddr) begin         // Hold low during write
      CCA_awready     <= #TCQ 1'b0;
    end else if (bsync_cfg_complete && !CCA_bvalid) begin // Release after write sync completes or write
      CCA_awready     <= #TCQ 1'b1;                       // response is accepted, whichever comes later.
    end
  end

  // Create wready output - hold low after data is captured until write completes
  // IP Checklist violation - Using unreg inputs (wvalid as part of wdata_active)
  always @(posedge cfg_clk) begin
    if (cfg_rst_q) begin
      CCA_wready      <= #TCQ 1'b0;
    end else if (set_ready_post_reset) begin              // Set to 1 after reset
      CCA_wready      <= #TCQ 1'b1;
    end else if (wdata_active || got_wdata) begin         // Hold low during write
      CCA_wready      <= #TCQ 1'b0;
    end else if (bsync_cfg_complete && !CCA_bvalid) begin // Release after write sync completes or write
      CCA_wready      <= #TCQ 1'b1;                       // response is accepted, whichever comes later.
    end
  end
  // }}} End Wait for Write Data/Address ---

  // {{{ Wait for Read Data ----------------
  // Start read sync process once address is available
  assign raddr_active = CF_arvalid && CCA_arready;
  assign rresp_active = CCA_rvalid  && CF_rready;

  // Capture read address from Config Fabric
  // No reset value necessary since read address not used until available
  //*ASSERTION*
  //(ap_raddr_sampled_incorrectly): cfg_raddr should be the same as the accepted address when sync_re asserts
  always @(posedge cfg_clk) begin
    if (CCA_arready) begin
      CCA_cfg_raddr   <= #TCQ {CF_araddr[23:2], 2'b0}; // Tying off lower bits results in less address decode logic
    end
  end

  // Create arready output - hold low after addr is captured until read completes
  // IP Checklist violation - Using unreg inputs (arvalid as part of raddr_active
  // and rready as part of rresp_active)
  //*ASSERTION*
  //(ap_arready_and_rvalid): rvalid is not asserted when arready is asserted
  // Note - this assertion precludes rresp_active AND raddr_active
  always @(posedge cfg_clk) begin
    if (cfg_rst_q) begin
      CCA_arready     <= #TCQ 1'b0;
    end else if (set_ready_post_reset) begin
      CCA_arready     <= #TCQ 1'b1;  // Set to 1 after reset
    end else if (raddr_active) begin // Clear when address received
      CCA_arready     <= #TCQ 1'b0;
    end else if (rresp_active) begin // Set when response transferred
      CCA_arready     <= #TCQ 1'b1;
    end
  end
  // }}} End Wait for Read Data ------------

  // {{{ Synchronization -------------------
  // {{{ + Write Sync + --------------------
  // {{{ ++ Write Data/Addr Sync ++ --------
  // Synchronize a read enable from the cfg_clk domain to the core_clk domain to know
  // when it's safe to sample the write address and data.

  // wsync_cfg_req asserts when the write address and data are accepted from the config
  // fabric. That signal is sampled in the core_clk domain and registered twice to
  // protect against metastability.  When the signal reaches the final core_clk domain
  // register stage (sync_we), the synchronizer is cleared. Since the signal asserts for
  // one core_clk cycle, it can be used directly as the write enable (indicating that the
  // write data and address have been stable long enough to sample them with core_clk).

  // Synchronize write enable to core_clk domain
  //*ASSERTION*
  //(ap_write_overlap): A new write is not received until the synchronization circuit is ready
  //(ap_lost_write_enable): sync_we is seen for every write
  always @(posedge cfg_clk or posedge CCA_sync_we) begin
    if (CCA_sync_we) begin
      wsync_cfg_req   <= #TCQ 1'b0;
    end else if (cfg_rst_q) begin             // cfg_rst_q will be put on D input b/c need async clr for synchronizer
      wsync_cfg_req   <= #TCQ 1'b0;
    end else if (set_we) begin
      wsync_cfg_req   <= #TCQ 1'b1;
    end
  end
  always @(posedge core_clk) begin
    if (CCA_sync_we) begin
      wsync_core_q    <= #TCQ 1'b0;
      CCA_sync_we     <= #TCQ 1'b0;
    end else begin
      wsync_core_q    <= #TCQ wsync_cfg_req;  // cfg_clk to core_clk domain crossing
      CCA_sync_we     <= #TCQ wsync_core_q;
    end
  end
  // }}} ++ End Write Data/Addr Sync ++ ----

  // {{{ ++ Write Ready Sync ++ ------------
  // We must not release the ready signals until the write is complete, so that the
  // address and data are held constant during the write.

  // bsync_cfg_req is a latched version of the synchronized write enable.
  // That signal is sampled in the cfg_clk domain and registered twice to protect against
  // metastability.  When the signal reaches the final cfg_clk domain register stage
  // (bsync_cfg_done), the synchronizer is cleared. We latch the resulting signal and use
  // it to indicate that the readys can be released (although that circuit also waits for
  // the config fabric to accept the write response).

  //*ASSERTION*
  //(ap_wready_overlap): A new write response is not initiated until the synchronization circuit is ready
  //(ap_lost_write_rdy_sync): A write ready release is seen for every sync_we
  always @(posedge core_clk or posedge bsync_cfg_done) begin
    if (bsync_cfg_done) begin
      bsync_core_req  <= #TCQ 1'b0;
    end else if (CCA_sync_cfg_rst) begin // CCA_sync_cfg_rst will be put on D input b/c need async clr for synchronizer
      bsync_core_req  <= #TCQ 1'b0;
    end else if (CCA_sync_we) begin
      bsync_core_req  <= #TCQ 1'b1;
    end
  end

  always @(posedge cfg_clk) begin
    if (bsync_cfg_done) begin
      bsync_cfg_q     <= #TCQ 1'b0;
      bsync_cfg_done  <= #TCQ 1'b0;
    end else begin
      bsync_cfg_q     <= #TCQ bsync_core_req;
      bsync_cfg_done  <= #TCQ bsync_cfg_q;
    end
  end

  always @(posedge cfg_clk) begin
    if (cfg_rst_q) begin
      bsync_cfg_hold_done <= #TCQ 1'b0;
    end else if (bsync_cfg_done) begin
      bsync_cfg_hold_done <= #TCQ 1'b1;
    end else if (bsync_cfg_hold_done && !CCA_bvalid) begin
      bsync_cfg_hold_done <= #TCQ 1'b0;
    end
  end

  assign bsync_cfg_complete = bsync_cfg_done || bsync_cfg_hold_done;
  // }}} ++ End Write Ready Sync ++ --------
  // }}} + End Write Sync + ----------------

  // {{{ + Read Sync+ ----------------------
  // Synchronize Config Fabric Read Interface - no relationship between
  // cfg_clk and core_clk is assumed.

  // {{{ ++ Read Address Sync ++ -----------
  // Synchronize a read enable from the cfg_clk domain to the core_clk domain to know
  // when it's safe to sample the read address.

  // arsync_cfg_req asserts when the read address is accepted from the config fabric.
  // That signal is sampled in the core_clk domain and registered twice to protect
  // against metastability.  When the signal reaches the final core_clk domain register
  // stage (sync_re), the synchronizer is cleared. Since the signal asserts for one
  // core_clk cycle, it can be used directly as the read enable (indicating that the read
  // address has been stable long enough for the read data to settle).

  //*ASSERTION*
  //(ap_read_overlap): A new read is not received until the synchronization circuit is ready
  //(ap_lost_read_enable): A sync_re is seen for every read
  always @(posedge cfg_clk or posedge CCA_sync_re) begin
    if (CCA_sync_re) begin
      arsync_cfg_req  <= #TCQ 1'b0;
    end else if (cfg_rst_q) begin     // cfg_rst_q will be put on D input b/c need async clr for synchronizer
      arsync_cfg_req  <= #TCQ 1'b0;
    end else if (raddr_active) begin
      arsync_cfg_req  <= #TCQ 1'b1;
    end
  end

  // Create read enable for read data assembly (check for rising edge of
  // synchronized read enable)
  always @(posedge core_clk) begin
    if (CCA_sync_re) begin            // Because of reset sync, it's ok to not reset these flops with CCA_sync_cfg_rst
      arsync_core_q   <= #TCQ 1'b0;   // (the writable reg bank will be held in reset long enough for sync to clear)
      CCA_sync_re     <= #TCQ 1'b0;
    end else begin
      arsync_core_q   <= #TCQ arsync_cfg_req;
      CCA_sync_re     <= #TCQ arsync_core_q;
   end
  end
  // }}} ++ End Read Address Sync ++ -------

  // {{{ ++ Read Response Sync ++ ----------
  // Synchronize the read enable back from the core_clk domain to the cfg_clk domain to
  // know when it's safe to sample the read data in order to form the read response.

  // rsync_cfg_req is a latched version of the synchronized read enable.
  // That signal is sampled in the cfg_clk domain and registered twice to protect against
  // metastability.  When the signal reaches the final cfg_clk domain register stage
  // (rsync_cfg_done), the synchronizer is cleared. Since the signal asserts for one
  // core_clk cycle, it can be used directly as the read enable (indicating that the read
  // address has been stable long enough for the read data to settle).

  //*ASSERTION*
  //(ap_rresp_overlap): A new read response is not initiated until the synchronization circuit is ready
  //(ap_lost_rresp): A read response sync done is seen for every sync_re
  always @(posedge core_clk or posedge rsync_cfg_done) begin
    if (rsync_cfg_done) begin                 // domain crossing
      rsync_core_req  <= #TCQ 1'b0;
    end else if (CCA_sync_cfg_rst) begin
      rsync_core_req  <= #TCQ 1'b0;
    end else if (CCA_sync_re) begin
      rsync_core_req  <= #TCQ 1'b1;
    end
  end

  // Synchronize read enable back to cfg_clk domain
  always @(posedge cfg_clk) begin
    if (rsync_cfg_done) begin
      rsync_cfg_q     <= #TCQ 1'b0;
      rsync_cfg_done  <= #TCQ 1'b0;
    end else begin
      rsync_cfg_q     <= #TCQ rsync_core_req; // domain crossing
      rsync_cfg_done  <= #TCQ rsync_cfg_q;
    end
  end
  // }}} ++ End Read Response Sync ++ ------
  // }}} + End Read Sync + -----------------
  // }}} End Synchronization ---------------

  // {{{ Write Response Generator ----------
  // Form write response with status OKAY when data and address are received.
  // Takes as input got_wdata and got_waddr.

  // Create bvalid output
  // Assert valid two cycles after data is received, clear on response transfer
  // IP Checklist violation - unreg input (bready) used
  //*COVERPOINT*
  //(cp_cf_backpressures_bresp): Config Fabric holds off write response by not immediately asserting ready
  //*ASSERTION*
  //(ap_resp_for_every_wdata): There is a write response for every write data received
  //(ap_resp_for_every_waddr): There is a write response for every write address received
  always @(posedge cfg_clk) begin
    if (cfg_rst_q) begin
      CCA_bvalid      <= #TCQ 1'b0;
    // Set when resp is synch'ed back to cfg_clk domain (only if readys are low in case rst happened mid-write)
    end else if (bsync_cfg_done && !CCA_awready && !CCA_wready && !cfg_rst_qq) begin
      CCA_bvalid      <= #TCQ 1'b1;
    end else if (CF_bready) begin
      CCA_bvalid      <= #TCQ 1'b0;
    end
  end
  // }}} End Write Response Generator ------

  // {{{ Read Response Generator -----------
  // Takes as input rsync_cfg_done (indicates when read data can safely be sampled)

  // Create rdata output
  // Get data from Read Data Assembly block. Safe to sample when rsync_cfg_done is
  // asserted.
  always @(posedge cfg_clk) begin
    if (cfg_rst_q) begin
      CCA_rdata       <= #TCQ 32'b0;
    // Refresh data when resp is synch'ed back to cfg_clk domain (only if ready is low in case rst happened mid-read)
    end else if (rsync_cfg_done && !CCA_arready && !cfg_rst_qq) begin
      CCA_rdata       <= #TCQ CC_core_rdata;
    end
  end

  // Create rvalid output when the read data is valid (rsync_cfg_done
  // asserts), clear on response transfer
  // IP Checklist violation - unreg input (rready) used
  //*COVERPOINT*
  //(cp_cf_backpressures_rresp): Config Fabric holds off response by not immediately asserting ready
  //*ASSERTION*
  //(ap_resp_for_every_read): There is a read response for every read
  always @(posedge cfg_clk) begin
    if (cfg_rst_q) begin
      CCA_rvalid      <= #TCQ 1'b0;
    // Set when resp is synch'ed back to cfg_clk domain (only if ready is low in case rst happened mid-read)
    end else if (rsync_cfg_done && !CCA_arready && !cfg_rst_qq) begin
      CCA_rvalid      <= #TCQ 1'b1;
    end else if (CF_rready) begin
      CCA_rvalid      <= #TCQ 1'b0;
    end
  end
  // }}} End Read Response Generator -------

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
//
// OLLM_RX_DATAPATH
// Description:
// This module holds most of the datapath functions and calculations
// for the OLLM_RX
//
// Hierarchy:
// PHY_TOP
//    |___OLLM_RX_TOP
//             |_____OLLM_RX_DATAPATH <-- this module
//             |_____OLLM_RX_ERR_DETECT
// ---------------------------------------------------------------------

`timescale 1ps/1ps

module srio_gen2_v4_1_16_ollm_rx_datapath
  #(
    parameter TCQ           = 100,  // in pS
    parameter IDLE1         = 1,    // Include the IDLE1 sequence {0, 1}
    parameter IDLE2         = 0,    // Include the IDLE2 sequence {0, 1}
    parameter VC            = 0,    // Highest number VC supported {0, 1}
    parameter SWITCH_MODE   = 0,    // If the core is generated with Switch Mode Support {0, 1}
    parameter RETRY         = 1,    // Includes Retry protocol {0, 1}
    parameter TARGET_DS     = 0,  
    parameter VC1_CT        = 1)    // Default traffic mode for VC1 {0, 1}
   (
  // {{{ port declarations ----------------
    // clocks and resets and general signals
    input             phy_clk,                    // PHY interface clock
    input             phy_rst_q,                  // Reset for PHY clock Domain
    output            PR_phy_rcvd_link_reset,     // Received 4 consecutive link reset control symbols
    output     [31:0] prd_debug,                  // OLLM RX Debug bus, should include useful signals for HW debug

    // OPLM/OLLM RX CS Decode Interface
    input      [63:0] PRD_rx_data,                // Receive data
    input      [7:0]  PRD_rx_charisk,             // Indicates which bytes are K characters
    input      [1:0]  PRD_rx_valid,               // Indicates valid words
    input      [81:0] PRD_cs_decode,              // A whole series of control symbol decodes. See assignment
    input             PRD_idle2_selected,         // Indicates when an IDLE2 sequence is present
    input             PP_out_of_sync,             // Scrambler is out of sync
    input             PP_port_initialized,        // Indicates port is initialized

    // RX Buffer Interface
    output reg        PR_phyr_tvalid,             // Valid data indicator
    input             BR_phyr_tready,             // Destination Ready
    output     [63:0] PR_phyr_tdata,              // Packet for transfer
    output reg [7:0]  PR_phyr_tkeep,              // Byte Enable for transferred packet
    output reg        PR_phyr_tlast,              // Last DW of incoming packet
    output reg [7:0]  PR_phyr_tuser,              // {1'h0, skip_crc, 3'h0, VC, CRF, src_dsc} AXI Compliance Pad
    input      [5:0]  BR_phy_buf_stat,            // Buffer status from the RX Buffer

    // OLLM TX Interface
    input             PT_sent_init_cs,            // Indicates we sent 15 control symbols
    output reg        PR_link_initialized,        // Indicates we are ready to transmit data
    output reg        PR_rewind,                  // An error or retry condition has been seen
    output reg [5:0]  PR_phy_rcvd_buf_stat,       // Buffer status received from the link partner
    output reg        PR_send_rfr,                // Send an RFR control symbol (Request)
    input             PT_rfr_sent,                // Sent RFR (Grant)
    output reg        PR_send_lreq,               // Send a Link Request Control Symbol
    input             PT_lreq_sent,               // Sent Link Request
    output reg        PR_send_pna,                // Send a PNA control symbol
    input             PT_pna_sent,                // Sent PNA
    output reg        PR_send_pr,                 // Send a PR control symbol
    input             PT_pr_sent,                 // Sent PR
    output reg        PR_send_lresp,              // Send a Link Response Control Symbol
    input             PT_lresp_sent,              // Sent Link Response
    output reg [4:0]  PR_port_stat,               // Current port status
    output reg        PR_port_stat_ok,            // Port status is specifically in the OK state
    output reg        PR_output_retry_stop,       // OLLM RX is currently in Output Retry Stopped State
    output reg        PR_output_error_stop,       // OLLM RX is currently in Output Error Stopped State
    output reg        PR_port_error,              // OLLM RX is currently in Port Error State
    output reg        PR_input_retry_stop,        // OLLM RX is currently in Input Retry Stopped State
    output reg        PR_input_error_stop,        // OLLM RX is currently in Input Error Stopped State
    output reg        PR_input_status_good,       // OLLM RX is currently in Input Waiting for Event State
    output reg        PR_rcvd_error_free_status,  // Asserts when an error free status control symbol is received

    // PHY Config Interface
    input             PC_load_ackids,             // Loads next_rcvd_pkt and last_ack with the CFG provided alternatives
    input             PC_clr_port_error,          // Clear the Output port error state
    input             PC_error_disable,           // Disable error checking in the OLLM RX
// FIXVC - next two signals currently unused
    input             PC_vc_ct,                   // VC1 is in continuous traffic mode and all VC1 should be acked
    input             PC_vc_en,                   // Enable VC1 operation
    output reg        PR_rcvd_lresp,              // Asserted when a link response has been received
    output reg [5:0]  PR_ackid_status,            // sampled from parameter0
    output reg [4:0]  PR_rcvd_port_stat,          // Last received link partner's port status
    output reg        PR_rcvd_pa_or_pna,          // Asserted when a Packet Accepted or Not Accepted has been received

    // internal connections to error detection block
    output     [1:0]  pd_flag_stg0,               // Packet Delimiter Delimiter indication
    output     [1:0]  sc_flag_stg0,               // Control Symbol Delimiter indication
    output     [1:0]  in_packet_stg0,             // Indicates when in or out of a packet
    output     [1:0]  sop,                        // successful decode of SOP in either upper or lower
    output     [1:0]  stomp,                      // successful decode of STOMP in either upper or lower
    output     [1:0]  eop,                        // successful decode of EOP in either upper or lower
    output     [1:0]  rfr,                        // successful decode of RFR in either upper or lower
    output     [1:0]  lreq,                       // successful decode of LREQ in either upper or lower
    output     [1:0]  stat,                       // successful decode of STAT in either upper or lower
    output     [1:0]  mce,                        // successful decode of MCE in either upper or lower
    // stage 1 inputs (packet CRC checking)
    output reg [63:0] masked_rx_data_stg1,        // Receive data, masked AckID for CRC check
    output reg [63:0] ordered_rx_data_stg1,       // Receive data
    output            data_vld_stg1,              // data valid window
    output reg [1:0]  data_vld_stg0_d,            // delayed data valid window to identify charisk
    output reg        data_stream_enable_stg1,    // stream enable for both RT and CT
    output reg        pp_out_of_sync_stg1,        // Scrambler is out of sync
    output reg        pp_port_initialized_stg1,   // Indicates port is initialized
    output reg [3:0]  crc_loc_stg1,               // one-hot location for the CRC
    output reg        mid_crc_loc_stg1,           // Beat identifier for the mid CRC
    output reg        beat_count_q_is_10,         // Just might be the location of the mid-crc
    output reg        framing_end_stg1,           // indicates the end of a packet
    output reg        framing_start_stg1,         // indicates the start of a packet
    output reg        framing_dsc_stg1,           // used with in_packet to indicate a discontinued packet
    output reg        upper_valid_stg1,           // Data valid signal after reordering for AXI
    output reg        lower_valid_stg1,           // Data valid signal after reordering for AXI
    output reg        lower_padded_stg1,          // when 1, the lower word is pad at the end of a packet
    output reg        first_beat_stg1,            // first beat of a packet
    output reg        stomp_detect_stg1,          // Stomp control symbol received
    output reg        lreq_detect_stg1,           // Link-Request detection
    output reg [1:0]  lreq_in_stat_detect_stg1,   // Link-Request detection - in stat
    output reg [1:0]  pa_detect_stg1,             // Packet-Ack identifier
    output     [1:0]  pa_detect_stg0,             // Packet-Ack identifier
    output reg        pr_detect_stg1,             // Packet-Retry identifier
    output reg        rfr_detect_stg1,            // Restart-from-Retry identifier
    output reg [5:0]  pa_ackid_stg1,              // sampled from parameter0 - pa ackid
    output reg [5:0]  pr_ackid_stg1,              // sampled from parameter0 - pr ackid
    output reg [1:0]  expected_ackid_coef_stg1,   // when two PAs, value of 2, otherwise 1
    // stage 2 inputs
    // stage 2
    output reg        lresp_detect_stg2,          // Link-Response identifier
    output reg        framing_end_stg2,           // used with in_packet to indicate the end of a packet
    output reg        framing_start_stg2,         // used with in_packet to indicate the start of a packet
    output reg  [3:0] crc_loc_stg2,               // one-hot location for the CRC
    output reg        mid_crc_loc_stg2,           // Beat identifier for the mid CRC
    output reg        rt_stream_enable_stg2,      // Used to enable the stream for RT
    output            dest_dsc_stg2,              // Determination for destination discontinue
    output reg        err_recovery,
    output reg        carryover_stg2,

    // outputs consumed by datapath
    input             prx_out_fatal_detect,       // Output fatal error condition discovered
    input             prx_force_send_lreq,        // Forces the OLLM TX to send a LREQ
    input             prx_out_recoverable_detect, // Output recoverable error condition discovered
    input             prx_in_recoverable_detect,  // Input recoverable error condition discovered
    input             prx_in_retry_detect,        // Retry condition discovered
    input       [3:0] prx_cs_crc_check_fail,      // used to generate cs_crc_in_error_cond
    input             prx_cs_in_error_cond,       // control symbol error condition detected
    input             prx_rcvd_bad_status,        // Asserts when there is an error in status
    output            in_retry_stopped_state,     // indicates the input error state as Retry Stopped
    input             idle2_sync_char_stg0,
    input             control_sym_in_error_cond_cmb,// This signal is asserted combo, when CS errors asserted
    output            not_in_retry_stopped_state,   // CR 825487, to check the next state of input error rec state machine
    input             idle_seq_in_error_cond_cmb,   // checks the idle seq errors combonatorally
    input             lreq_pd_error,                // this signal detects the PD erros in LREQ
    output      [1:0] lreq_reset_dev,               // LREQ + RST condition detection
    output            in_error_stopped_state,       // added to fix the CR# 837481
    input             idle2_7_4_beat_err_cmb        //
  // }}} ----------------------------------
   );

  // {{{ local parameters -----------------

  // Special Character decodes
  localparam [7:0] PD                    = 8'b011_11100; // K28.3
  localparam [7:0] SC                    = 8'b000_11100; // K28.0
  localparam [7:0] K_CHAR                = 8'b101_11100; // K28.5
  localparam [7:0] R_CHAR                = 8'b111_11101; // K29.7
  localparam [7:0] A_CHAR                = 8'b111_11011; // K27.7
  localparam [7:0] M_CHAR                = 8'b001_11100; // K28.1

  // Stype1 decodes
  localparam [2:0] C_SOP                 = 3'b000;
  localparam [2:0] C_STMP                = 3'b001;
  localparam [2:0] C_EOP                 = 3'b010;
  localparam [2:0] C_RFR                 = 3'b011;
  localparam [2:0] C_LREQ                = 3'b100;
  localparam [2:0] C_MCE                 = 3'b101;
  localparam [2:0] C_RSVD1               = 3'b110;
  localparam [2:0] C_NOP                 = 3'b111;

  // Stype0 decodes
  localparam [2:0] C_PA                  = 3'b000;
  localparam [2:0] C_PR                  = 3'b001;
  localparam [2:0] C_PNA                 = 3'b010;
  localparam [2:0] C_RSVD0               = 3'b011;
  localparam [2:0] C_STAT                = 3'b100;
  localparam [2:0] C_VSTAT               = 3'b101;
  localparam [2:0] C_LRESP               = 3'b110;
  localparam [2:0] C_IMP_DEF             = 3'b111;

  // CMD decodes
  localparam [2:0] C_LREQ_RST_DEV        = 3'b011; // sub-command for link request
  localparam [2:0] C_LREQ_IN_STAT        = 3'b100; // sub-command for link request

  // Output Error Handler States
  localparam [5:0] OUT_RECOVERY_DISABLED = 6'b000001;
  localparam [5:0] OUT_WAIT_FOR_EVENT    = 6'b000010;
  localparam [5:0] OUT_STOP_ERROR        = 6'b000100;
  localparam [5:0] OUT_ERROR_RECOVER     = 6'b001000;
  localparam [5:0] OUT_STOP_RETRY        = 6'b010000;
  localparam [5:0] OUT_FATAL             = 6'b100000;

  // Input Error Handler States
  localparam [6:0] IN_RECOVERY_DISABLED  = 7'b0000001;
  localparam [6:0] IN_WAIT_FOR_EVENT     = 7'b0000010;
  localparam [6:0] IN_STOP_INPUT         = 7'b0000100;
  localparam [6:0] IN_ERROR_STOPPED      = 7'b0001000;
  localparam [6:0] IN_ERROR_RECOVERY     = 7'b0010000;
  localparam [6:0] IN_RETRY_STOPPED      = 7'b0100000;
  localparam [6:0] IN_REC_DISABLED_LRESP = 7'b1000000;

  // Port Status
  localparam [4:0] PORT_STAT_ERROR       = 5'b00010;
  localparam [4:0] PORT_STAT_RETRY_STOP  = 5'b00100;
  localparam [4:0] PORT_STAT_ERROR_STOP  = 5'b00101;
  localparam [4:0] PORT_STAT_OK          = 5'b10000;

  // FTYPE Decode
  localparam [3:0] NREAD                 = 4'b0010;
  localparam [3:0] NWRITE                = 4'b0101;
  localparam [3:0] SWRITE                = 4'b0110;
  localparam [3:0] MAINTENANCE           = 4'b1000;
  localparam [3:0] DSTREAM               = 4'b1001;
  localparam [3:0] DOORBELL              = 4'b1010;
  localparam [3:0] MESSAGE               = 4'b1011;
  localparam [3:0] RESPONSE              = 4'b1101;


  // }}} End local parameters -------------


  // {{{ wire declarations ----------------
  // Prefix notation:
  // phy   = phy clock domain
  // pr/PR = Physical Layer Receive
  // pt/PT = Physical Layer Transmit
  // pc/PC = Physical Layer Config
  // pp/PP = Physical Layer OPLM
  // br/BR = Buffer Layer Receive
  // prx   = Physical Layer Error Detection signals (Not 'pre' to avoid confusion)
  // _stg* = Pipeline Stage Number

  // Pipeline stage 0 signals
  //wire  [1:0]            pd_flag_stg0;             // Packet Delimiter Delimiter indication
  //wire  [1:0]            sc_flag_stg0;             // Control Symbol Delimiter indication

  // - Stype1 Decode
  //wire  [1:0]            in_packet_stg0;           // indicates when the the data stream is part of a packet
  wire                   framing_start_stg0;       // used with in_packet to indicate the start of a packet
  wire                   framing_end_stg0;         // used with in_packet to indicate the end of a packet
  wire                   framing_dsc_stg0;         // used with in_packet to indicate a discontinued packet
  wire                   framing_dsc_stg0_delay;   // used with in_packet to indicate a discontinued packet
  wire  [1:0]            data_vld_stg0;            // data valid window, based off of in_packet
  //wire  [1:0]            sop;                     // successful decode of SOP in either upper or lower
  //wire  [1:0]            stomp;                   // successful decode of STOMP in either upper or lower
  //wire  [1:0]            eop;                     // successful decode of EOP in either upper or lower
  //wire  [1:0]            rfr;                     // successful decode of RFR in either upper or lower
  //wire  [1:0]            lreq;                    // successful decode of LREQ in either upper or lower
  wire  [1:0]            lreq_rst_dev;             // successful decode of LREQ-rst-dev in either upper or lower
  wire  [1:0]            lreq_in_stat;             // successful decode of LREQ-in-stat in either upper or lower
  //wire  [1:0]            mce;                      // successful decode of MCE in either upper or lower
  wire  [1:0]            s1rsvd;                   // successful decode of RSVD in either upper or lower
  wire  [1:0]            nop;                      // successful decode of NOP in either upper or lower

  // - Stype0 Decode
  wire  [5:0]            pa_ackid_stg0;            // sampled from parameter0 - pa ackid
  wire  [5:0]            pr_ackid_stg0;            // sampled from parameter0 - pr ackid
  wire  [5:0]            ackid_status_stg0;        // sampled from parameter0
  wire  [2:0]            vcid_stg0;                // sampled from parameter0
  wire  [4:0]            port_status_stg0;         // sampled from parameter1
  wire  [5:0]            buf_status_stg0;          // sampled from parameter1
  wire  [4:0]            cause_stg0;               // sampled from parameter1
  wire  [1:0]            pa;                       // successful decode of PA in either upper or lower
  wire  [1:0]            pr;                       // successful decode of PR in either upper or lower
  wire  [1:0]            pna;                      // successful decode of PNA in either upper or lower
  wire  [1:0]            s0rsvd;                   // successful decode of RSVD in either upper or lower
  //wire  [1:0]            stat;                    // successful decode of STATUS in either upper or lower
  wire  [1:0]            vcstat;                   // successful decode of VC STATUS in either upper or lower
  wire  [1:0]            lresp;                    // successful decode of LRESP in either upper or lower
  wire  [1:0]            id;                       // successful decode of ID in either upper or lower
  wire                   standard_dsc_case;//CR 821476

  // - Link Initialization
  reg   [2:0]            rcvd_good_status_cnt;     // counter used to determine if link initialization is complete
  reg   [2:0]            rcvd_good_status_cnt_q;   // counter used to determine if link initialization is complete


  // Pipeline stage 1 signals
  // - Carryover from Stage 0
  reg   [1:0]            pd_flag_stg1;             // Packet Delimiter Delimiter indication
  //reg                    pp_out_of_sync_stg1;      // Scrambler is out of sync
  //reg                    pp_port_initialized_stg1; // Indicates port is initialized
  reg                    enable_state_stg1;        // Tells the input state machine to stay in its current state

  reg   [1:0]            in_packet_stg1;           // indicates when the the data stream is part of a packet
  //reg                    framing_start_stg1;       // used with in_packet to indicate the start of a packet
  //reg                    framing_end_stg1;         // used with in_packet to indicate the end of a packet
  //reg                    framing_dsc_stg1;         // used with in_packet to indicate a discontinued packet
  //reg   [5:0]            pa_ackid_stg1;            // sampled from parameter0 - pa ackid
  //reg   [5:0]            pr_ackid_stg1;            // sampled from parameter0 - pr ackid
  reg   [2:0]            vcid_stg1;                // sampled from parameter0
  reg   [5:0]            buf_status_stg1;          // sampled from parameter1
  reg                    update_buf_stat_stg1;     // indicates when it's ok to update
  reg   [4:0]            cause_stg1;               // sampled from parameter1
  reg   [4:0]            port_status_stg1;         // sampled from parameter1
  reg   [1:0]            lresp_detect_stg1;        // Link-Response detection
  //reg                    lreq_detect_stg1;         // Link-Request detection - in stat
  //reg   [1:0]            lreq_in_stat_detect_stg1; // Link-Request detection
  //reg                    rfr_detect_stg1;          // RFR detection
  reg                    pna_detect_stg1;          // PNA detection
  //reg                    pr_detect_stg1;           // PR detection
  reg   [1:0]            pr_detect_lanes_stg1;     // PR detection
  //reg   [1:0]            pa_detect_stg1;           // PA detection
  //reg                    stomp_detect_stg1;        // PA detection
  //reg                    mid_crc_loc_stg1;         // Beat identifier for the mid CRC

  // - Data Formatter
  //reg   [3:0]            crc_loc_stg1;             // one-hot location for the CRC
  reg                    user_def_stg1;            // signal indicates a user defined packet
  reg  [31:0]            carryover_data_stg1;      // Storage for an extra Word
  reg                    carryover_stg1;           // Indicates if carryover_data is fresh or stale
  //reg                    upper_valid_stg1;         // Data valid signal after reordering for AXI
  //reg                    lower_valid_stg1;         // Data valid signal after reordering for AXI
  //reg                    lower_padded_stg1;        // when 1, the lower word is pad at the end of a packet
  //reg                    first_beat_stg1;          // first beat of a packet
  reg                    first_beat_stg1_early;    // first beat of a packet
  //reg  [63:0]            ordered_rx_data_stg1;     // Receive data, reordered for AXI
  //reg  [63:0]            masked_rx_data_stg1;      // Receive data, reordered for AXI, masked AckID for CRC check
  reg                    eop_partial_stg1;         // End-of-Packet, incomplete
  reg                    dsc_partial_stg1;         // Packet Discontinue, incomplete
//  reg                    data_stream_enable_stg1;  // stream enable for both RT and CT
  reg                    vc_stg1;                  // VC, pulled from data stream
  reg                    crf_stg1;                 // CRF, pulled from data stream
  wire                   qualified_data_vld_stg1;  // combined data_vld signal - at least one word is valid
  reg                    single_cycle_stg1;        // When asserted, only one beat of data will go out on AXI
  reg                    first_beat_stg1_d;        // Find the first beat of a packet
  reg                    first_beat_stg1_early_d;  // Find the first beat of a packet
//  reg                    standard_dsc_case_delay;//CR 821476
  reg                    prx_in_recoverable_detect_delay  ;//CR 821476

  // Pipeline stage 2 signals
  // - Carryover from Stage 1
  reg                    in_packet_stg2;           // indicates when the the data stream is part of a packet
  reg  [63:0]            ordered_rx_data_stg2;     // Receive data, reordered for AXI
//  reg   [3:0]            crc_loc_stg2;             // one-hot location for the CRC
  reg                    user_def_stg2;            // signal indicates a user defined packet
  reg                    data_vld_stg2;            // combined data_vld signal - at least one word is valid
  //reg                    framing_start_stg2;       // used with in_packet to indicate the start of a packet
  //reg                    framing_end_stg2;         // used with in_packet to indicate the end of a packet
  reg                    framing_dsc_stg2;         // used with in_packet to indicate a discontinued packet
  reg                    framing_dsc_stg3;         // used with in_packet to indicate a discontinued packet
  reg   [5:0]            buf_status_stg2;          // sampled from parameter1
  reg   [4:0]            cause_stg2;               // sampled from parameter1
  reg                    lreq_in_stat_detect_stg2; // Link-Request detection
  reg                    lreq_in_stat_detect_stg2_bit0; // Link-Request detection // new signal
  reg                    lreq_in_stat_detect_stg2_bit1; // Link-Request detection // new signal
//  reg                    carryover_stg2;           // Indicates if carryover_data is fresh or stale
  reg                    lower_padded_stg2;        // when 1, the lower word is pad at the end of a packet
  reg                    lower_padded_stg2_spec;   // speculative - when 1, the lower word is pad at the end of a packet
  reg                    set_eop_stg2;             // complete End-of-Packet determination
  reg                    eop_delay_stg2;           // delay eop by one cycle
  reg                    set_dsc_stg2;             // discontinue due to stomp, lreq, rfr
  reg                    dsc_delay_stg2;           // delay dsc by one cycle
  reg                    vc_stg2;                  // VC, pulled from data stream
  reg                    crf_stg2;                 // CRF, pulled from data stream
  //reg                    mid_crc_loc_stg2;         // Beat identifier for the mid CRC
  reg                    single_cycle_stg2;        // When asserted, only one beat of data will go out on AXI
  reg                    first_beat_stg2;          // first beat of a packet
  reg                    pr_detect_stg2;           // PR detection
  reg   [1:0]            pr_detect_lanes_stg2;     // PR detection
  reg                    pna_detect_stg2;          // PNA detection
  //reg                    lresp_detect_stg2;        // Link-Response detection

  // - Input Error Handler - FSM
  //reg                    rt_stream_enable_stg2;    // Used to enable the stream for RT

  // Pipeline stage 3 signals
  // - Carryover from Stage 2
  reg                    in_packet_stg3;           // indicates when the the data stream is part of a packet
  reg  [63:0]            ordered_rx_data_stg3;     // Receive data, reordered for AXI
  reg   [3:0]            crc_loc_stg3;             // one-hot location for the CRC
  reg                    data_vld_stg3;            // combined data_vld signal - at least one word is valid
  reg                    framing_start_stg3;       // used with in_packet to indicate the start of a packet
  reg                    framing_end_stg3;         // used with in_packet to indicate the end of a packet
  reg                    lower_padded_stg3;        // when 1, the lower word is pad at the end of a packet
  reg                    set_eop_stg3;             // complete End-of-Packet determination
  reg                    eop_delay_stg3;           // delay eop by one cycle
  reg                    set_dsc_stg3;             // discontinue due to stomp, lreq, rfr
  reg                    vc_stg3;                  // VC, pulled from data stream
  reg                    crf_stg3;                 // CRF, pulled from data stream
  reg                    dest_dsc_stg3;            // Determination for destination discontinue
  reg                    mid_crc_loc_stg3;         // Beat identifier for the mid CRC
  reg                    single_cycle_stg3;        // When asserted, only one beat of data will go out on AXI
  reg                    rt_stream_enable_stg3;    // Used to enable the stream for RT
  reg                    large_packet_stg3;        // Asserts when a packet exceeds 80 bytes
  reg                    lresp_detect_stg3;        // Link-Response detection
  reg   [1:0]            pr_detect_lanes_stg3;     // PR detection

  // Pipeline stage 4 signals

  // - RX Buf Interface
  reg   [3:0]            crc_loc_stg4;             // one-hot location for the CRC
  reg                    large_packet_stg4;        // Asserts when a packet exceeds 80 bytes
  reg  [63:0]            phyr_tdata;               // un-swizzled data going to the buffer
  reg                    pr_phyr_tlast_d;          // combinatorial version of TLAST
  wire                   advance_condition;        // circumstance by which the AXI bus should advance
  reg                    out_of_packet;            // indicates when not in a packet on the buffer interface
  reg  [1:0]             eop_q;
  // }}} End wire declarations ------------


  // {{{ prd_debug assignment --------------
  assign prd_debug = {24'h0,
                      PR_input_retry_stop,
                      PR_input_error_stop,
                      PR_output_retry_stop,
                      PR_output_error_stop,
                      pr_detect_stg2,
                      PR_send_pr,
                      pna_detect_stg2,
                      PR_send_pna};

  // }}} -----------------------------------


// {{{ Stage0 Pipeline -------------------

  // {{{ + CS Decode Demux ------------------

  assign pd_flag_stg0        = PRD_cs_decode[81:80];
  assign sc_flag_stg0        = PRD_cs_decode[79:78];

  assign in_packet_stg0      = PRD_cs_decode[77:76];
  assign framing_start_stg0  = PRD_cs_decode[75];
  assign framing_end_stg0    = PRD_cs_decode[74];
  assign framing_dsc_stg0    = PRD_cs_decode[73];
  assign sop                 = PRD_cs_decode[72:71];
  assign stomp               = PRD_cs_decode[70:69];
  assign eop                 = PRD_cs_decode[68:67];
  assign rfr                 = PRD_cs_decode[66:65];
  assign lreq                = PRD_cs_decode[64:63];
  assign lreq_rst_dev        = PRD_cs_decode[62:61];
  assign lreq_reset_dev      = PRD_cs_decode[62:61];//
  assign lreq_in_stat        = PRD_cs_decode[60:59];
  assign mce                 = PRD_cs_decode[58:57];
  assign s1rsvd              = PRD_cs_decode[56:55];
  assign nop                 = PRD_cs_decode[54:53];

  assign pa_ackid_stg0       = PRD_cs_decode[52:47];
  assign pr_ackid_stg0       = PRD_cs_decode[46:41];
  assign ackid_status_stg0   = PRD_cs_decode[40:35];
  assign vcid_stg0           = PRD_cs_decode[34:32];
  assign port_status_stg0    = PRD_cs_decode[31:27];
  assign buf_status_stg0     = PRD_cs_decode[26:21];
  assign cause_stg0          = PRD_cs_decode[20:16];
  assign pa                  = PRD_cs_decode[15:14] & {2{PR_link_initialized}};
  assign pr                  = PRD_cs_decode[13:12] & {2{PR_link_initialized}};
  assign pna                 = PRD_cs_decode[11:10] & {2{PR_link_initialized}};
  assign s0rsvd              = PRD_cs_decode[9:8];
  assign stat                = PRD_cs_decode[7:6];
  assign vcstat              = PRD_cs_decode[5:4];
  assign lresp               = PRD_cs_decode[3:2];
  assign id                  = PRD_cs_decode[1:0];

  // STYPE1 Coverage:

    // *- COVERAGE (cp_PR_short_stype1_in_upper)
    // Observe every type of short control symbol in upper

    // *- COVERAGE (cp_PR_short_stype1_in_lower)
    // Observe every type of short control symbol in lower

    // *- COVERAGE (cp_PR_long_stype1_in_upper)
    // Observe every type of long control symbol starting in upper

    // *- COVERAGE (cp_PR_long_stype1_in_lower)
    // Observe every type of long control symbol starting in lower

    // *- COVERAGE (cp_PR_cross_short_stype1_upper_lower)
    // Observe two short control symbol in both positions, cross all types

    // *- COVERAGE (cp_PR_cross_short_stype1_consecutive)
    // Observe a short control symbol in lower, followed by short control
    // symbol in upper of next data beat, cross all types

    // *- COVERAGE (cp_PR_lreq_as_eop)
    // Observe lreq (in-stat and reset-dev) as a packet delimiter in both IDLE1 and IDLE2
    // both in and out of input error state

    // *- coverage (cp_pr_rfr_as_eop)
    // observe rfr as a packet delimiter in both IDLE1 and IDLE2
    // both in and out of input retry state

    // *- coverage (cp_pr_stomp_as_eop)
    // observe stomp as a packet delimiter in both IDLE1 and IDLE2
    // both in and out of input retry state

    // *- COVERAGE (cp_PR_cs_after_sop_1)
    // Observe sop control symbol followed by one non packet delimiting control symbol

    // *- COVERAGE (cp_PR_cs_after_sop_2)
    // Observe sop control symbol followed by two non packet delimiting control symbols

    // *- COVERAGE (cp_PR_cs_after_sop_3)
    // Observe sop control symbol followed by three non packet delimiting control symbols

    // *- COVERAGE (cp_PR_cs_after_sop_4)
    // Observe sop control symbol followed by four non packet delimiting control symbols

    // *- COVERAGE (cp_PR_cs_before_eop_1)
    // Observe eop control symbol preceded by one non packet delimiting control symbol

    // *- COVERAGE (cp_PR_cs_before_eop_2)
    // Observe eop control symbol preceded by two non packet delimiting control symbols

    // *- COVERAGE (cp_PR_cs_before_eop_3)
    // Observe eop control symbol preceded by three non packet delimiting control symbols

    // *- COVERAGE (cp_PR_cs_before_eop_4)
    // Observe eop control symbol preceded by four non packet delimiting control symbols

    // *- COVERAGE (cp_PR_cs_before_sop_1)
    // Observe sop, used to end a packet and start a new packet, preceded by one non packet delimiting control symbols

    // *- COVERAGE (cp_PR_cs_before_sop_2)
    // Observe sop, used to end a packet and start a new packet, preceded by two non packet delimiting control symbols

    // *- COVERAGE (cp_PR_cs_before_sop_3)
    // Observe sop, used to end a packet and start a new packet, preceded by three non packet delimiting control symbols

    // *- COVERAGE (cp_PR_cs_before_sop_4)
    // Observe sop, used to end a packet and start a new packet, preceded by four non packet delimiting control symbols

    // *- COVERAGE (cp_PR_cs_mid_packet_upper)
    // Observe a non packet delimiting control symbol in the middle of framed data in the upper half

    // *- COVERAGE (cp_PR_cs_mid_packet_lower)
    // Observe a non packet delimiting control symbol in the middle of framed data in the lower half

    // *- COVERAGE (cp_PR_cs_out_of_packet_upper)
    // Observe a non packetdelimiting control symbol outside of framed data in the upper half

    // *- COVERAGE (cp_PR_cs_out_of_packet_lower)
    // Observe a non packet delimiting control symbol outside of framed data in the lower half

    // *- COVERAGE (cp_PR_cs_after_1_data)
    // Observe one word of data after sof, followed by a non packet delimiting control symbol

    // *- COVERAGE (cp_PR_cs_after_2_data)
    // Observe two words of data after sof, followed by a non packet delimiting control symbol

    // *- COVERAGE (cp_PR_cs_before_1_data)
    // Observe a non packet control symbol followed by one word of data, followed by an end delimiter

    // *- COVERAGE (cp_PR_cs_before_2_data)
    // Observe a non packet control symbol followed by two words of data, followed by an end delimiter

    // *- COVERAGE (cp_PR_reset_device_scenario1)
    // Observe four consecutive Link-Request reset-device control symbols

    // *- COVERAGE (cp_PR_reset_device_scenario2)
    // Observe four Link-Request reset-device control symbols, separated by status/NOP control symbols

    // *- COVERAGE (cp_PR_reset_device_scenario3)
    // Observe four Link-Request reset-device control symbols, seperated by other control symbols control symbols

    // *- COVERAGE (cp_PR_start_and_end)
    // Observe framing_start_stg0 and framing_end_stg0 on the same cycle

    // *- COVERAGE (cp_PR_start_1before_end)
    // Observe framing_start_stg0 one cycle before framing_end_stg0

    // *- COVERAGE (cp_PR_start_2before_end)
    // Observe framing_start_stg0 two cycle before framing_end_stg0

    // *- COVERAGE (cp_PR_start_1after_end)
    // Observe framing_start_stg0 one cycle after framing_end_stg0

    // *- COVERAGE (cp_PR_start_2after_end)
    // Observe framing_start_stg0 two cycle after framing_end_stg0


  // STYPE0 Coverage:

    // *- COVERAGE (cp_PR_short_stype0_in_upper)
    // Observe every type of short control symbol in upper

    // *- COVERAGE (cp_PR_short_stype0_in_lower)
    // Observe every type of short control symbol in lower

    // *- COVERAGE (cp_PR_long_stype0_in_upper)
    // Observe every type of long control symbol starting in upper

    // *- COVERAGE (cp_PR_long_stype0_in_lower)
    // Observe every type of long control symbol starting in lower

    // *- COVERAGE (cp_PR_cross_short_stype0_upper_lower)
    // Observe two short control symbols in both positions, cross all types

    // *- COVERAGE (cp_PR_cross_short_stype0_consecutive)
    // Observe a short control symbol in lower, followed by short control
    // symbol in upper of next data beat, cross all types

    // *- COVERAGE (cp_PR_stype1_in_packet)
    // Observe every type of control symbol while in-packet

    // *- COVERAGE (cp_PR_stype1_out_of_packet)
    // Observe every type of control symbol while out-of-packet


  // }}} End of CS Decode Demux -----------


  // {{{ + Data Valid Generation ------------

  // Data Valid - When in packet, mask out any inter-packet control symbols
  assign data_vld_stg0 = {in_packet_stg0[1] && !PRD_rx_charisk[7] && !PRD_rx_charisk[4],
                          in_packet_stg0[0] && !PRD_rx_charisk[3] && !PRD_rx_charisk[0]};

  // }}} End of Data Valid Generation -----


  // {{{ + Link Reset Detection -------------

  // by specification, we must see four consecutive LREQ-reset-device
  // control symbols in order to qualify a true reset-device request.
  // Any other symbols interwoven in the four causes the count to be cleared.
  reg [2:0] reset_device_cnt;

  assign PR_phy_rcvd_link_reset = reset_device_cnt[2];
  wire clear_rst_cnt0 = (pd_flag_stg0[0] || sc_flag_stg0[0]) && (!(stat[0] && nop[0]) && !lreq_rst_dev[0]);
  wire clear_rst_cnt1 = (pd_flag_stg0[1] || sc_flag_stg0[1]) && (!(stat[1] && nop[1]) && !lreq_rst_dev[1]);
  always @(posedge phy_clk) begin
    if (phy_rst_q)
      reset_device_cnt <= #TCQ 3'b000;
    else if (!PR_link_initialized)
      reset_device_cnt <= #TCQ 3'b000;
    // special case - clear condition in upper and reset req in lower, clear previous and reload with 1 (for lower)
    else if (clear_rst_cnt1 && lreq_rst_dev[0])
      reset_device_cnt <= #TCQ 3'b001;
    else if (clear_rst_cnt1)
      reset_device_cnt <= #TCQ 3'b000;
    // special case - if there's a clear condition in the lower only clear if the upper isn't the 4th reset
    else if (clear_rst_cnt0 && !(lreq_rst_dev[1] && reset_device_cnt == 3'h3))
      reset_device_cnt <= #TCQ 3'b000;
    else if (&lreq_rst_dev)
      reset_device_cnt <= #TCQ {1'b0, reset_device_cnt[1:0]} + 2;
    else if (|lreq_rst_dev)
      reset_device_cnt <= #TCQ {1'b0, reset_device_cnt[1:0]} + 1;
    else if (PR_phy_rcvd_link_reset)
      reset_device_cnt <= #TCQ {1'b0, reset_device_cnt[1:0]};
  end

  // }}} End of Link Reset Detection ------


  // {{{ + Link Initialization --------------

  always @(posedge phy_clk) begin
    if (phy_rst_q)
      PR_link_initialized <= #TCQ 1'b0;
    else if (!PP_port_initialized)
      PR_link_initialized <= #TCQ 1'b0;
    else if (PT_sent_init_cs && (rcvd_good_status_cnt == 3'h7) && !prx_rcvd_bad_status)
      PR_link_initialized <= #TCQ 1'b1;
  end

  reg stat_q, stat_qq;
  reg prx_rcvd_bad_status_q, prx_rcvd_bad_status_qq;
  reg pr_rcvd_error_free_status_d;
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      stat_q                    <= #TCQ 1'b0;
      stat_qq                   <= #TCQ 1'b0;
      prx_rcvd_bad_status_q     <= #TCQ 1'b0;
      prx_rcvd_bad_status_qq    <= #TCQ 1'b0;
      PR_rcvd_error_free_status <= #TCQ 1'b0;
      rcvd_good_status_cnt_q    <= #TCQ 3'h0;
    end else begin
      stat_q                    <= #TCQ |stat;
      stat_qq                   <= #TCQ stat_q;
      prx_rcvd_bad_status_q     <= #TCQ prx_rcvd_bad_status;
      prx_rcvd_bad_status_qq    <= #TCQ prx_rcvd_bad_status_q;
      PR_rcvd_error_free_status <= #TCQ pr_rcvd_error_free_status_d && !prx_rcvd_bad_status;
      rcvd_good_status_cnt_q    <= #TCQ rcvd_good_status_cnt;
    end
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      rcvd_good_status_cnt        <= #TCQ 3'h0;
      pr_rcvd_error_free_status_d <= #TCQ 1'b0;
    end else if (!PP_port_initialized) begin
      rcvd_good_status_cnt        <= #TCQ 3'h0;
      pr_rcvd_error_free_status_d <= #TCQ 1'b0;
    end else if (rcvd_good_status_cnt_q != 3'h7 &&
                 (prx_cs_in_error_cond || prx_rcvd_bad_status || prx_rcvd_bad_status_qq)) begin
      rcvd_good_status_cnt        <= #TCQ 3'h0;
      pr_rcvd_error_free_status_d <= #TCQ 1'b0;
    end else if (stat_qq && rcvd_good_status_cnt != 3'h7 && !prx_in_recoverable_detect) begin
      rcvd_good_status_cnt        <= #TCQ rcvd_good_status_cnt + 1;
      pr_rcvd_error_free_status_d <= #TCQ 1'b1;
    end else if (rcvd_good_status_cnt_q != 3'h7 && prx_in_recoverable_detect) begin
      rcvd_good_status_cnt        <= #TCQ 3'h0;
    end else begin
      pr_rcvd_error_free_status_d <= #TCQ 1'b0;
    end
  end


    // *- COVERAGE (cp_PR_link_initialization_sequence)
    // Observe a proper link initialization sequence

    // *- COVERAGE (cp_PR_link_initialization_error_sequence)
    // Observe an error condition crossed with rcvd_good_status = {0, 1, 2, 6, 7}

    // *- COVERAGE (cp_PR_port_initialization_dropped)
    // Observe PP_port_intialized drop crossed with rcvd_good_status = {0, 1, 2, 6, 7}

    // *- COVERAGE (cp_PR_link_reinitialization)
    // Observe reinitialization after PP_port_intialized reasserts

    // *- COVERAGE (cp_PR_link_initialization_b2b)
    // Observe back to back status on link initialization


  // }}} End of Link Initialization -------

// }}} End Stage0 Pipeline ---------------


// {{{ Stage1 Pipeline -------------------

  // {{{ + Stage1 Pipeline Registers --------
  // register the inputs to the OPLM interface.
  always @(posedge phy_clk) begin
    pp_out_of_sync_stg1         <= #TCQ PP_out_of_sync;
    pp_port_initialized_stg1    <= #TCQ PP_port_initialized;
  end

  // register signals created by stage 0 logic.
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      pd_flag_stg1              <= #TCQ 2'h0;
      in_packet_stg1            <= #TCQ 2'h0;
      framing_start_stg1        <= #TCQ 1'b0;
      framing_end_stg1          <= #TCQ 1'b0;
      framing_dsc_stg1          <= #TCQ 1'b0;
      pa_ackid_stg1             <= #TCQ 6'h3F;
      pr_ackid_stg1             <= #TCQ 6'h3F;
      PR_ackid_status           <= #TCQ 6'h00;
      update_buf_stat_stg1      <= #TCQ 1'b0;
      vcid_stg1                 <= #TCQ 3'h0;
      cause_stg1                <= #TCQ 5'h00;
      port_status_stg1          <= #TCQ 5'h10;
      PR_rcvd_port_stat         <= #TCQ 5'h10;
      lresp_detect_stg1         <= #TCQ 2'h0;
      PR_rcvd_lresp             <= #TCQ 1'b0;
      lreq_detect_stg1          <= #TCQ 1'b0;
      lreq_in_stat_detect_stg1  <= #TCQ 2'h0;
      rfr_detect_stg1           <= #TCQ 1'b0;
      pna_detect_stg1           <= #TCQ 1'b0;
      pr_detect_stg1            <= #TCQ 1'b0;
      pr_detect_lanes_stg1      <= #TCQ 2'h0;
      pa_detect_stg1            <= #TCQ 2'h0;
      stomp_detect_stg1         <= #TCQ 1'b0;
      expected_ackid_coef_stg1  <= #TCQ 2'h0;
      enable_state_stg1         <= #TCQ 1'b0;
      eop_q                     <= #TCQ 2'h0;
      data_vld_stg0_d           <= #TCQ 2'h0;
    end else begin

      pd_flag_stg1              <= #TCQ pd_flag_stg0;

      // from stype1 decode
      in_packet_stg1            <= #TCQ in_packet_stg0;
      framing_start_stg1        <= #TCQ framing_start_stg0;
      framing_end_stg1          <= #TCQ framing_end_stg0 && data_stream_enable_stg1;
      framing_dsc_stg1          <= #TCQ framing_dsc_stg0 && data_stream_enable_stg1;

      // from stype0 decode
      pa_ackid_stg1             <= #TCQ pa_ackid_stg0;
      pr_ackid_stg1             <= #TCQ pr_ackid_stg0;
      PR_ackid_status           <= #TCQ ackid_status_stg0;
      vcid_stg1                 <= #TCQ vcid_stg0;
      update_buf_stat_stg1      <= #TCQ (|pa || |pr || |stat);
      cause_stg1                <= #TCQ cause_stg0;
      port_status_stg1          <= #TCQ port_status_stg0;
      PR_rcvd_port_stat         <= #TCQ port_status_stg0;
      // Added !(PRD_idle2_selected && PP_out_of_sync) to fix the CR# 838891
      // All control symbols and packet received while a lane descrambler in IDLE2 is
      // out of sync shall be ignored and discarded. Spec 6, 4.8.3 //
      lresp_detect_stg1         <= #TCQ lresp & {2{!(PRD_idle2_selected && pp_out_of_sync_stg1)}};//
      PR_rcvd_lresp             <= #TCQ |lresp && PR_link_initialized;
      lreq_detect_stg1          <= #TCQ |lreq & {2{!(PRD_idle2_selected && pp_out_of_sync_stg1)}};//
      lreq_in_stat_detect_stg1  <= #TCQ lreq_in_stat;
      rfr_detect_stg1           <= #TCQ |rfr & {2{!(PRD_idle2_selected && pp_out_of_sync_stg1)}};//
      pna_detect_stg1           <= #TCQ |pna & {2{!(PRD_idle2_selected && pp_out_of_sync_stg1)}};//
      pr_detect_stg1            <= #TCQ |pr & {2{!(PRD_idle2_selected && pp_out_of_sync_stg1)}};//
      pr_detect_lanes_stg1      <= #TCQ pr;
     // pa_detect_stg1            <= #TCQ pa & {2{!(PRD_idle2_selected && pp_out_of_sync_stg1)}};//12/18/2014
      pa_detect_stg1            <= #TCQ pa & {2{!(PRD_idle2_selected && (PP_out_of_sync || pp_out_of_sync_stg1))}};
      stomp_detect_stg1         <= #TCQ |stomp & {2{!(PRD_idle2_selected && pp_out_of_sync_stg1)}};//
      expected_ackid_coef_stg1  <= #TCQ &pa ? 2'h2 : 2'h1;
      enable_state_stg1         <= #TCQ PR_link_initialized;
      eop_q                     <= #TCQ eop;
      data_vld_stg0_d           <= #TCQ data_vld_stg0;
    end
  end

  assign pa_detect_stg0 = pa & {2{!(PRD_idle2_selected && pp_out_of_sync_stg1)}};//

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      buf_status_stg1 <= #TCQ 6'h00;
    end else if (|pa || |pr || |stat) begin
      buf_status_stg1 <= #TCQ buf_status_stg0;
    end else if (|prx_cs_crc_check_fail[2:0] || prx_cs_in_error_cond) begin
      buf_status_stg1 <= #TCQ buf_status_stg2;
    end else if (prx_cs_crc_check_fail[3]) begin
      buf_status_stg1 <= #TCQ PR_phy_rcvd_buf_stat;
    end
  end


  // }}} End of Stage1 Pipeline Registers -
  // Added below code as part of CR# 842999 fix. The idle2_sync_char_stg0 appears
  // only in IDLE2 condition.
  reg idle2_sync_char_stg1;
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
        idle2_sync_char_stg1 <= 1'b0;
    end else begin
        idle2_sync_char_stg1 <= idle2_sync_char_stg0;
    end
  end
  // {{{ + Data Formatter -------------------

  // Generate the carryover logic -
  // These are shadow registers used to hold extra data when
  // building packet data to go to the buffer. There are scenarios
  // where we can have three words when we only have enough bandwidth
  // for two. In these cases, we store the extra word until the next cycle.
  // Two scenarios exist for having carryover data.
  always @(posedge phy_clk) begin
    carryover_data_stg1    <= #TCQ PRD_rx_data[31:0];
    if (phy_rst_q) begin
      carryover_stg1 <= #TCQ 1'b0;
    // cases under which we may have to store more than two meaningful words
    // scenario 1. We are already in a carryover state
    // scenario 2. One valid word is stored, waiting for another word
    end else if (!data_stream_enable_stg1) begin
      carryover_stg1 <= #TCQ 1'b0;
    // added to fix the CR# 842999, when sync sequence is detected in IDLE2, the packet is cancelled
    // so there is no need to store any data beats
    // no need to add protection of PRD_idle2_selected as idle2_sync_char_stg0 is generated only in IDLE2.
    end else if (idle2_sync_char_stg1) begin
      carryover_stg1 <= #TCQ 1'b0;
    end else if (carryover_stg1 || (upper_valid_stg1 && !lower_valid_stg1)) begin
      // a. Two valid pieces of data arrive OR
      // b. Observe end of a packet/start of a new packet (via solo SOP)
      //     and a valid word arrives for the beginning of the next packet
      if (&data_vld_stg0 || (framing_end_stg0 && data_vld_stg0[0])) begin
        carryover_stg1 <= #TCQ 1'b1;
      end else begin
        carryover_stg1 <= #TCQ 1'b0;
      end
    end
  end

  wire stomp_pulse;

  assign stomp_pulse = |stomp && !stomp_detect_stg1;

  reg stomp_pulse_stg1;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
        stomp_pulse_stg1 <= #TCQ 1'b0;
    end else begin
        stomp_pulse_stg1 <= #TCQ stomp_pulse;
    end
  end

  // organize the phy data -
  // Pack everything from MSB to LSB.
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      upper_valid_stg1     <= #TCQ 1'b0;
      lower_valid_stg1     <= #TCQ 1'b0;
      ordered_rx_data_stg1 <= #TCQ 64'h0;
      masked_rx_data_stg1  <= #TCQ 64'h0;
      lower_padded_stg1    <= #TCQ 1'b0;
      vc_stg1              <= #TCQ 1'b0;
      crf_stg1             <= #TCQ 1'b0;

    //end else if ((!data_stream_enable_stg1 && !framing_start_stg0)) begin
    //added (PRD_idle2_selected && |lreq) condition to discard the valid stage in IDLE2 cases //
    //added lreq_detect_stg1 || stomp_detect_stg1 to fix CR 825747
    end else if ((!data_stream_enable_stg1 && !framing_start_stg0)
                 ||
                 //lreq_detect_stg1 || stomp_detect_stg1 // <-- replaced this logic with below line //
                 (lreq[1] && !PRD_idle2_selected) ||   // fix for CR 842990
                 (lreq[0] && !carryover_stg1 && !PRD_idle2_selected) ||
                 (stomp_pulse_stg1 && !PRD_idle2_selected)
                 ||
                 (PRD_idle2_selected && (|lreq) && !carryover_stg1)//
                 //(PRD_idle2_selected && |lreq)//
                 ) begin
      upper_valid_stg1     <= #TCQ 1'b0;
      lower_valid_stg1     <= #TCQ 1'b0;
      lower_padded_stg1    <= #TCQ 1'b0;

    // if there is a carryover, it automatically goes in the upper location
    // The lower location will hold the next piece of valid data from stage1
    end else if (carryover_stg1) begin
      ordered_rx_data_stg1[63:32]  <= #TCQ carryover_data_stg1;
      masked_rx_data_stg1[63:32]   <= #TCQ first_beat_stg1_d ?
                                           {6'h00, carryover_data_stg1[25:0]} : carryover_data_stg1;
      upper_valid_stg1             <= #TCQ 1'b1;
      vc_stg1                      <= #TCQ 1'b0; // first_beat_stg1_d ? carryover_data_stg1[25] && (VC == 1) : vc_stg1;
      crf_stg1                     <= #TCQ first_beat_stg1_d ? carryover_data_stg1[24] : crf_stg1;
      if (data_vld_stg0[1]) begin
        ordered_rx_data_stg1[31:0] <= #TCQ PRD_rx_data[63:32];
        masked_rx_data_stg1[31:0]  <= #TCQ PRD_rx_data[63:32];
        lower_valid_stg1           <= #TCQ 1'b1;
        lower_padded_stg1          <= #TCQ 1'b0;
      // pad last word, use stale data
      // looking for framing_end_stg0 without the extra overhead
      end else if ((in_packet_stg0[1] && pd_flag_stg0[1]) || (in_packet_stg0[0] && pd_flag_stg0[0])) begin
        lower_valid_stg1           <= #TCQ 1'b1;
        lower_padded_stg1          <= #TCQ 1'b1;
        if (in_packet_stg0[1] && pd_flag_stg0[1])             // CR 806709
        ordered_rx_data_stg1[31:0] <= #TCQ PRD_rx_data[63:32];// CR 806709
        if (in_packet_stg0[0] && pd_flag_stg0[0])                 // CR 806709
        ordered_rx_data_stg1[31:0] <= #TCQ PRD_rx_data[31:0]; // CR 806709

      end else if (data_vld_stg0[0]) begin
        ordered_rx_data_stg1[31:0] <= #TCQ PRD_rx_data[31:0];
        masked_rx_data_stg1[31:0]  <= #TCQ PRD_rx_data[31:0];
        lower_valid_stg1           <= #TCQ 1'b1;
        lower_padded_stg1          <= #TCQ 1'b0;
      end else begin
        lower_valid_stg1           <= #TCQ 1'b0;
        lower_padded_stg1          <= #TCQ 1'b0;
      end

    // if we currently are holding one valid piece of data in stage2 -
    // find the next piece of valid data from stage1 and store it in lower
    end else if (upper_valid_stg1 && !lower_valid_stg1) begin
      if (data_vld_stg0[1]) begin
        ordered_rx_data_stg1[31:0] <= #TCQ PRD_rx_data[63:32];
        masked_rx_data_stg1[31:0]  <= #TCQ PRD_rx_data[63:32];
        lower_valid_stg1           <= #TCQ 1'b1;
        lower_padded_stg1          <= #TCQ 1'b0;
      // pad last word, use stale data
      // looking for framing_end_stg0 without the extra overhead
      end else if ((in_packet_stg0[1] && pd_flag_stg0[1]) || (in_packet_stg0[0] && pd_flag_stg0[0])) begin
        lower_valid_stg1           <= #TCQ 1'b1;
        lower_padded_stg1          <= #TCQ 1'b1;
        if (in_packet_stg0[1] && pd_flag_stg0[1])             // CR 806709
        ordered_rx_data_stg1[31:0] <= #TCQ PRD_rx_data[63:32];// CR 806709
        if (in_packet_stg0[0] && pd_flag_stg0[0])                 // CR 806709
        ordered_rx_data_stg1[31:0] <= #TCQ PRD_rx_data[31:0]; // CR 806709

      end else if (data_vld_stg0[0]) begin
        ordered_rx_data_stg1[31:0] <= #TCQ PRD_rx_data[31:0];
        masked_rx_data_stg1[31:0]  <= #TCQ PRD_rx_data[31:0];
        lower_valid_stg1           <= #TCQ 1'b1;
        lower_padded_stg1          <= #TCQ 1'b0;
      end else begin
        lower_valid_stg1           <= #TCQ 1'b0;
        lower_padded_stg1          <= #TCQ 1'b0;
      end

    // if both upper and lower stage2 valids are 1 or 0 (treated the same) -
    // fill upper first, followed by lower
    end else begin
      if (data_vld_stg0[1]) begin
        ordered_rx_data_stg1[63:32] <= #TCQ PRD_rx_data[63:32];
        ordered_rx_data_stg1[31:0]  <= #TCQ PRD_rx_data[31:0];
        masked_rx_data_stg1[63:32]  <= #TCQ first_beat_stg1_d ? {6'h00, PRD_rx_data[57:32]} : PRD_rx_data[63:32];
        vc_stg1                     <= #TCQ first_beat_stg1_d ? PRD_rx_data[57] && (VC == 1) : vc_stg1;
        crf_stg1                    <= #TCQ first_beat_stg1_d ? PRD_rx_data[56] : crf_stg1;
        upper_valid_stg1            <= #TCQ PRD_idle2_selected ? !(|lreq) : 1'b1;//!idle2_sync_char_stg0;//1'b1;//!(|lreq);//
        masked_rx_data_stg1[31:0]   <= #TCQ PRD_rx_data[31:0];
        lower_valid_stg1            <= #TCQ data_vld_stg0[0] || pd_flag_stg0[0];
        lower_padded_stg1           <= #TCQ pd_flag_stg0[0];
      end else if (data_vld_stg0[0]) begin
        ordered_rx_data_stg1[63:32] <= #TCQ PRD_rx_data[31:0];
        masked_rx_data_stg1[63:32]  <= #TCQ (first_beat_stg1_d || pd_flag_stg0[1]) ?
                                             {6'h00, PRD_rx_data[25:0]} : PRD_rx_data[31:0];
        vc_stg1                     <= #TCQ (first_beat_stg1_d || pd_flag_stg0[1]) ?
                                             PRD_rx_data[25] && (VC == 1) : vc_stg1;
        crf_stg1                    <= #TCQ (first_beat_stg1_d || pd_flag_stg0[1]) ? PRD_rx_data[24] : crf_stg1;
        upper_valid_stg1            <= #TCQ 1'b1;
        lower_valid_stg1            <= #TCQ 1'b0;
        lower_padded_stg1           <= #TCQ 1'b0;
      end else if (!(lower_valid_stg1 && !data_vld_stg1)) begin
        upper_valid_stg1            <= #TCQ 1'b0;
        lower_valid_stg1            <= #TCQ 1'b0;
        lower_padded_stg1           <= #TCQ 1'b0;
      end
    end
  end


  // Partial generation of EOP -
  // Generation of the EOP straddles over two pipeline stages
  // because an EOP can arrive many cycles after the actual last
  // piece of data, with which it is associated. If EOP arrives
  // from the OPLM and this logic is still bundling up the last
  // DWORD of data, this section handles it. If the last piece of
  // data has already been bundled, we have to forward EOP to the
  // next cycle
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      eop_partial_stg1 <= #TCQ 1'b0;
      dsc_partial_stg1 <= #TCQ 1'b0;
    end else if (carryover_stg1) begin
      eop_partial_stg1 <= #TCQ framing_end_stg0 && data_stream_enable_stg1;
      dsc_partial_stg1 <= #TCQ framing_dsc_stg0;
    end else if (upper_valid_stg1 && !qualified_data_vld_stg1) begin
      eop_partial_stg1 <= #TCQ framing_end_stg0 && data_stream_enable_stg1;
      dsc_partial_stg1 <= #TCQ framing_dsc_stg0;
    end else if (data_vld_stg0[1]) begin
      eop_partial_stg1 <= #TCQ framing_end_stg0 && data_stream_enable_stg1;
      dsc_partial_stg1 <= #TCQ framing_dsc_stg0;
    end else begin
      eop_partial_stg1 <= #TCQ 1'b0;
    end
  end


  // turn of the data valid when in an error or recovery state, or when
  // not initialized yet. This also depends on what VC mode is running in
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      data_stream_enable_stg1 <= #TCQ 1'b0;
    end else if (!rt_stream_enable_stg2) begin
      data_stream_enable_stg1 <= #TCQ 1'b0;
    end else if (framing_start_stg0) begin
      // FIXVC - add PC value to see if in CT
      if (vc_stg1) begin
        data_stream_enable_stg1 <= #TCQ PR_link_initialized;
      end else begin
        data_stream_enable_stg1 <= #TCQ rt_stream_enable_stg2;
      end
    end
  end

  // wait to push data out until we have collected two words AND
  // we are certain that the EOP doesn't need to advance.
  // You can do that by waiting for at least one more word of data to arrive.
  //
  // This is a very timing-sensitive signal. The logic here is not what would be
  // usually used if we didn't have such a tough timing path.
  wire embedded_control_symbols  = // set when there are control symbols in both the upper and lower
                             (PRD_rx_charisk[7] && (PRD_rx_charisk[3] || PRD_idle2_selected)) ||
                             (PRD_rx_charisk[4] && PRD_rx_charisk[3] && PRD_idle2_selected);
  assign data_vld_stg1           = lower_valid_stg1 && // upper_valid is 1 when lower_valid is 1
                             (!embedded_control_symbols || carryover_stg1 || framing_end_stg1 ||
                             (!carryover_stg1 && PRD_rx_charisk[7] && |pd_flag_stg0));
  assign qualified_data_vld_stg1 = data_stream_enable_stg1 && data_vld_stg1;


  // find the first beat of a packet so we can grab stream details
  always @* begin
    if (framing_end_stg0 && !carryover_stg1 && data_vld_stg0[0] &&
        !(upper_valid_stg1 && !lower_valid_stg1) && !first_beat_stg1) begin
      first_beat_stg1_d       = 1'b1;
      first_beat_stg1_early_d = 1'b1;
    end else if ((framing_end_stg1 || (framing_end_stg0 && !data_stream_enable_stg1)) &&
                 !first_beat_stg1_early) begin
      first_beat_stg1_d       = 1'b1;
      first_beat_stg1_early_d = 1'b0;
    end else if (qualified_data_vld_stg1) begin
      first_beat_stg1_d       = 1'b0;
      first_beat_stg1_early_d = 1'b0;
    end else begin
      first_beat_stg1_d       = first_beat_stg1;
      first_beat_stg1_early_d = 1'b0;
    end
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      first_beat_stg1       <= #TCQ 1'b1;
      first_beat_stg1_early <= #TCQ 1'b1;
    end else begin
      first_beat_stg1       <= #TCQ first_beat_stg1_d;
      first_beat_stg1_early <= #TCQ first_beat_stg1_early_d;
    end
  end

    // *- COVERAGE (cp_PR_carryover_asserts_one_cycle)
    // Observe that the carryover signal is asserted for one data beat

    // *- COVERAGE (cp_PR_carryover_asserts_multi_cycle)
    // Observe that the carryover signal is asserted for more than one data beat

    // *- COVERAGE (cp_PR_carryover_cross_data_vld)
    // Cross carryover_stg1 with data_vld_stg0 and framing_end_stg0

    // *- COVERAGE (cp_PR_carryover_before_lower_padded)
    // Observe carryover_stg1 asserted one cycle before lower_padded_stg1

    // *- COVERAGE (cp_PR_not_carryover_before_lower_padded)
    // Observe that carryover_stg1 is not asserted one cycle before lower_padded_stg1


  // }}} End of Data Formatter ------------


  reg  [4:0] beat_count, beat_count_q;
  wire [3:0] ftype_stg1 = ordered_rx_data_stg1[51:48];
  wire       tt_stg1    = ordered_rx_data_stg1[52];
  wire [3:0] ttype_stg1 = tt_stg1 ? ordered_rx_data_stg1[15:12] : ordered_rx_data_stg1[31:28];
  generate if (TARGET_DS == 1) begin: data_streaming_on
  // {{{ + CRC Location Finder --------------

  // CRC location finder -
  // There can be 32 bits of padding in either the upper or lower
  // as well as 16 bits of padding in either the first or third quadrant.
  // There are three conditions which determine the location of the
  // CRC within the DWORD: FTYPE, TT[0], and if packet size is >80 bytes
  // FTYPE = 2/8,   TT[0] = 0,     : crc_loc = 0100
  // FTYPE = 2/8,   TT[0] = 1,     : crc_loc = 0010
  // FTYPE = 5,     TT[0] = 0, <80 : crc_loc = 0100
  // FTYPE = 5,     TT[0] = 0, >80 : crc_loc = 0010
  // FTYPE = 5,     TT[0] = 1, <80 : crc_loc = 0010
  // FTYPE = 5,     TT[0] = 1, >80 : crc_loc = 0001
  // FTYPE = 6,     TT[0] = 0, <80 : crc_loc = 1000
  // FTYPE = 6,     TT[0] = 0, >80 : crc_loc = 0100
  // FTYPE = 6,     TT[0] = 1, <80 : crc_loc = 0100
  // FTYPE = 6,     TT[0] = 1, >80 : crc_loc = 0010
  // FTYPE = 10,    TT[0] = 0,     : crc_loc = 1000
  // FTYPE = 10,    TT[0] = 1,     : crc_loc = 0100
  // FTYPE = 11/13, TT[0] = 0, <80 : crc_loc = 0001
  // FTYPE = 11/13, TT[0] = 0, >80 : crc_loc = 1000
  // FTYPE = 11/13, TT[0] = 1, <80 : crc_loc = 1000
  // FTYPE = 11/13, TT[0] = 0, >80 : crc_loc = 0100
  reg  [5:0] crc_loc_logic, crc_loc_logic_q; 
  wire [1:0] start_end = tt_stg1 ? ordered_rx_data_stg1[7:6] : ordered_rx_data_stg1[23:22];
  wire       odd_stg1 = tt_stg1 ? ordered_rx_data_stg1[1] : ordered_rx_data_stg1[17];

  always @* begin
    if (first_beat_stg1 && lower_valid_stg1 && data_stream_enable_stg1) begin
      casex ({ftype_stg1, tt_stg1,odd_stg1,start_end})
      {NREAD, 1'b0, 1'bx, 2'bxx}       : crc_loc_logic = 6'b00_0100;
      {NREAD, 1'b1, 1'bx, 2'bxx}       : crc_loc_logic = 6'b00_0010;

      {NWRITE, 1'b0, 1'bx, 2'bxx}      : crc_loc_logic = 6'b00_0100;
      {NWRITE, 1'b1, 1'bx, 2'bxx}      : crc_loc_logic = 6'b00_0010;

      {SWRITE, 1'b0, 1'bx, 2'bxx}      : crc_loc_logic = 6'b00_1000;
      {SWRITE, 1'b1, 1'bx, 2'bxx}      : crc_loc_logic = 6'b00_0100;

      {DSTREAM, 1'b0, 1'b0, 2'b00}      : crc_loc_logic = 6'b10_0000; // Data stream & 8-bit devID
      {DSTREAM, 1'b0, 1'b0, 2'b01}      : crc_loc_logic = 6'b10_0001; // Data stream & 8-bit devID
      {DSTREAM, 1'b0, 1'b0, 2'b1x}      : crc_loc_logic = 6'b10_0010; // Data stream & 8-bit devID
      {DSTREAM, 1'b0, 1'b1, 2'b00}      : crc_loc_logic = 6'b10_0100; // Data stream & 8-bit devID
      {DSTREAM, 1'b0, 1'b1, 2'b01}      : crc_loc_logic = 6'b10_0101; // Data stream & 8-bit devID
      {DSTREAM, 1'b0, 1'b1, 2'b1x}      : crc_loc_logic = 6'b10_0110; // Data stream & 8-bit devID

      {DSTREAM, 1'b1, 1'b0, 2'b00}      : crc_loc_logic = 6'b10_1000; // Data stream & 16-bit devID
      {DSTREAM, 1'b1, 1'b0, 2'b01}      : crc_loc_logic = 6'b10_1001; // Data stream & 16-bit devID
      {DSTREAM, 1'b1, 1'b0, 2'b1x}      : crc_loc_logic = 6'b10_1010; // Data stream & 16-bit devID
      {DSTREAM, 1'b1, 1'b1, 2'b00}      : crc_loc_logic = 6'b10_1100; // Data stream & 16-bit devID
      {DSTREAM, 1'b1, 1'b1, 2'b01}      : crc_loc_logic = 6'b10_1101; // Data stream & 16-bit devID
      {DSTREAM, 1'b1, 1'b1, 2'b1x}      : crc_loc_logic = 6'b10_1110; // Data stream & 16-bit devID

      {MAINTENANCE, 1'b0, 1'bx, 2'bxx}  : crc_loc_logic = 6'b00_0100;
      {MAINTENANCE, 1'b1, 1'bx, 2'bxx}  : crc_loc_logic = 6'b00_0010;

      {DOORBELL, 1'b0, 1'bx, 2'bxx}     : crc_loc_logic = 6'b00_1000;
      {DOORBELL, 1'b1, 1'bx, 2'bxx}     : crc_loc_logic = 6'b00_0100;

      {MESSAGE, 1'b0, 1'bx, 2'bxx}      : crc_loc_logic = 6'b00_0001;
      {MESSAGE, 1'b1, 1'bx, 2'bxx}      : crc_loc_logic = 6'b00_1000;

      {RESPONSE, 1'b0, 1'bx, 2'bxx}     : crc_loc_logic = 6'b00_0001;
      {RESPONSE, 1'b1, 1'bx, 2'bxx}     : crc_loc_logic = 6'b00_1000;


      // user defined - go and find the crc (that's why the upper bit is set)
      default             : crc_loc_logic = 6'b01_0001;
      endcase
    end else if (beat_count == 5'd10 && !beat_count_q_is_10 && !crc_loc_logic_q[4] && !crc_loc_logic_q[5]) begin
      crc_loc_logic = {crc_loc_logic_q[5:4], crc_loc_logic_q[0], crc_loc_logic_q[3:1]};
    end else begin
      crc_loc_logic = crc_loc_logic_q;
    end
  end


  always @(posedge phy_clk) begin
    if (phy_rst_q)
      crc_loc_logic_q <= #TCQ 6'b01_0001;
    else if (!vc_stg2 && !rt_stream_enable_stg2)
      crc_loc_logic_q <= #TCQ 6'b00_0001;
    else begin
        crc_loc_logic_q <= #TCQ crc_loc_logic;
    end
end

wire crc_pad;

assign crc_pad = ((crc_loc_logic == 6'b10_0100) || (crc_loc_logic == 6'b10_0010) ||
                 (crc_loc_logic == 6'b10_0001) || (crc_loc_logic == 6'b10_1000) ||
                 (crc_loc_logic == 6'b10_1110) || (crc_loc_logic == 6'b10_1101));

reg final_crc_pad;   	   
reg final_crc_pad_q;   	   

 always @(posedge phy_clk) begin
    if (phy_rst_q)
      final_crc_pad_q <= #TCQ 1'b0;
    else 
      final_crc_pad_q <= #TCQ final_crc_pad;
 end



  always @* begin
    if (first_beat_stg1 && lower_valid_stg1 && data_stream_enable_stg1) 
       final_crc_pad =  crc_pad;
    else if (beat_count_q == 5'd10) 
       final_crc_pad =  ~crc_pad;
     else
       final_crc_pad =  final_crc_pad_q;
     end

  always @* begin
    // user defined scenario. We assume crc to be in either the 0 or 2 position,
    // depending of if there is pad or not.
    if (crc_loc_logic_q[4] && !crc_loc_logic_q[5]) begin // This is the user-def bit
      if (lower_padded_stg1) begin
        crc_loc_stg1  = {crc_loc_logic_q[1:0], crc_loc_logic_q[3:2]};
        user_def_stg1 = crc_loc_logic_q[4];
      end else begin
        crc_loc_stg1  = crc_loc_logic_q[3:0]; // always 4'b0001
        user_def_stg1 = crc_loc_logic_q[4];
      end
    end else begin

 if (crc_loc_logic_q[5]) begin // This is the ftype9 bit
      if (lower_padded_stg1) begin
	 if (final_crc_pad)
             crc_loc_stg1  = 4'b1000;
	 else 
             crc_loc_stg1  = 4'b0100;

      end else begin
	 if (final_crc_pad)
             crc_loc_stg1  = 4'b0010;
	 else 
             crc_loc_stg1  = 4'b0001;
      end
    end

      else begin 
      crc_loc_stg1  = crc_loc_logic_q[3:0]; 
      user_def_stg1 = 1'b0;
     end
   end
 end
 end endgenerate //data streaming on ends



 generate if (TARGET_DS == 0) begin: data_streaming_off
  // {{{ + CRC Location Finder --------------

  // CRC location finder -
  // There can be 32 bits of padding in either the upper or lower
  // as well as 16 bits of padding in either the first or third quadrant.
  // There are three conditions which determine the location of the
  // CRC within the DWORD: FTYPE, TT[0], and if packet size is >80 bytes
  // FTYPE = 2/8,   TT[0] = 0,     : crc_loc = 0100
  // FTYPE = 2/8,   TT[0] = 1,     : crc_loc = 0010
  // FTYPE = 5,     TT[0] = 0, <80 : crc_loc = 0100
  // FTYPE = 5,     TT[0] = 0, >80 : crc_loc = 0010
  // FTYPE = 5,     TT[0] = 1, <80 : crc_loc = 0010
  // FTYPE = 5,     TT[0] = 1, >80 : crc_loc = 0001
  // FTYPE = 6,     TT[0] = 0, <80 : crc_loc = 1000
  // FTYPE = 6,     TT[0] = 0, >80 : crc_loc = 0100
  // FTYPE = 6,     TT[0] = 1, <80 : crc_loc = 0100
  // FTYPE = 6,     TT[0] = 1, >80 : crc_loc = 0010
  // FTYPE = 10,    TT[0] = 0,     : crc_loc = 1000
  // FTYPE = 10,    TT[0] = 1,     : crc_loc = 0100
  // FTYPE = 11/13, TT[0] = 0, <80 : crc_loc = 0001
  // FTYPE = 11/13, TT[0] = 0, >80 : crc_loc = 1000
  // FTYPE = 11/13, TT[0] = 1, <80 : crc_loc = 1000
  // FTYPE = 11/13, TT[0] = 0, >80 : crc_loc = 0100
  reg  [4:0] crc_loc_logic, crc_loc_logic_q; // upper bit used for user def crc detection
  always @* begin
    if (first_beat_stg1 && lower_valid_stg1 && data_stream_enable_stg1) begin
      case ({ftype_stg1, tt_stg1})
      {NREAD, 1'b0}       : crc_loc_logic = 5'b0_0100;
      {NREAD, 1'b1}       : crc_loc_logic = 5'b0_0010;

      {NWRITE, 1'b0}      : crc_loc_logic = 5'b0_0100;
      {NWRITE, 1'b1}      : crc_loc_logic = 5'b0_0010;

      {SWRITE, 1'b0}      : crc_loc_logic = 5'b0_1000;
      {SWRITE, 1'b1}      : crc_loc_logic = 5'b0_0100;

      {MAINTENANCE, 1'b0} : crc_loc_logic = 5'b0_0100;
      {MAINTENANCE, 1'b1} : crc_loc_logic = 5'b0_0010;

      {DOORBELL, 1'b0}    : crc_loc_logic = 5'b0_1000;
      {DOORBELL, 1'b1}    : crc_loc_logic = 5'b0_0100;

      {MESSAGE, 1'b0}     : crc_loc_logic = 5'b0_0001;
      {MESSAGE, 1'b1}     : crc_loc_logic = 5'b0_1000;

      {RESPONSE, 1'b0}    : crc_loc_logic = 5'b0_0001;
      {RESPONSE, 1'b1}    : crc_loc_logic = 5'b0_1000;

      // user defined - go and find the crc (that's why the upper bit is set)
      default             : crc_loc_logic = 5'b1_0001;
      endcase
    end else if (beat_count == 5'd10 && !beat_count_q_is_10 && !crc_loc_logic_q[4]) begin
      crc_loc_logic = {1'b0, crc_loc_logic_q[0], crc_loc_logic_q[3:1]};
    end else begin
      crc_loc_logic = crc_loc_logic_q;
    end
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q)
      crc_loc_logic_q <= #TCQ 5'b1_0001;
    else if (!vc_stg2 && !rt_stream_enable_stg2)
      crc_loc_logic_q <= #TCQ 5'b0_0001;
    else
      crc_loc_logic_q <= #TCQ crc_loc_logic;
  end


  always @* begin
    // user defined scenario. We assume crc to be in either the 0 or 2 position,
    // depending of if there is pad or not.
    if (crc_loc_logic_q[4]) begin // This is the user-def bit
      if (lower_padded_stg1) begin
        crc_loc_stg1  = {crc_loc_logic_q[1:0], crc_loc_logic_q[3:2]};
        user_def_stg1 = crc_loc_logic_q[4];
      end else begin
        crc_loc_stg1  = crc_loc_logic_q[3:0]; // always 4'b0001
        user_def_stg1 = crc_loc_logic_q[4];
      end
    end else begin
      crc_loc_stg1  = crc_loc_logic_q[3:0];
      user_def_stg1 = 1'b0;
    end
  end
 end endgenerate //data streaming off ends

  // count the beats until we find the mid-CRC - always the 81st and 82nd byte
  always @(*) begin
    if (framing_start_stg1 && (!qualified_data_vld_stg1 || framing_end_stg1)) begin
      beat_count       = 5'h0;
      mid_crc_loc_stg1 = qualified_data_vld_stg1 && beat_count_q_is_10;
    end else if (!PR_port_stat_ok) begin
      beat_count       = 5'h0;
      mid_crc_loc_stg1 = 1'b0;
    end else if (framing_start_stg1 && qualified_data_vld_stg1) begin
      beat_count       = 5'h1;
      mid_crc_loc_stg1 = 1'b0;
    end else if (qualified_data_vld_stg1) begin
      beat_count       = beat_count_q + 1;
      mid_crc_loc_stg1 = beat_count_q_is_10;
    end else begin
      beat_count       = beat_count_q;
      mid_crc_loc_stg1 = mid_crc_loc_stg2;
    end
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      beat_count_q               <= #TCQ 0;
      beat_count_q_is_10         <= #TCQ 1'b0;
    end else begin
      beat_count_q               <= #TCQ beat_count;
      beat_count_q_is_10         <= #TCQ beat_count == 5'd10;
    end
  end


  // single beat transfer -
  // Identify when there is only going to be a single beat for a transfer to the buffer.
  // Need to delay single-beat transfers in order to properly find the crc.
  // Single cycle transfers:
  // Response with no data
  always @(*) begin
    if (first_beat_stg1 && lower_valid_stg1 && data_stream_enable_stg1) begin
      single_cycle_stg1 = ((ftype_stg1 == RESPONSE) && (ttype_stg1 == 4'h0)) ||
                          ((ftype_stg1 == DOORBELL) && !tt_stg1) ||
                           framing_end_stg1;
    end else if (ftype_stg1 != RESPONSE) begin
      single_cycle_stg1 = 1'b0;
    end else begin
      single_cycle_stg1 = single_cycle_stg2;
    end
  end


  // }}} End of CRC Location Finder -------

// }}} End Stage1 Pipeline ---------------

wire input_error_state;

// {{{ Stage2 Pipeline -------------------

  // {{{ + Stage2 Pipeline Registers --------

  // register signals created by stage 0 logic.
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PR_rcvd_pa_or_pna        <= #TCQ 1'b0;
      data_vld_stg2            <= #TCQ 1'b0;
      in_packet_stg2           <= #TCQ 1'b0;
      framing_start_stg2       <= #TCQ 1'b0;
      framing_end_stg2         <= #TCQ 1'b0;
      framing_dsc_stg2         <= #TCQ 1'b0;
      framing_dsc_stg3         <= #TCQ 1'b0;// new signal RC fix
      cause_stg2               <= #TCQ 5'h00;
      lreq_in_stat_detect_stg2 <= #TCQ 1'b0;
      PR_phy_rcvd_buf_stat     <= #TCQ 6'h0;
      user_def_stg2            <= #TCQ 1'b0;
      carryover_stg2           <= #TCQ 1'b0;
      mid_crc_loc_stg2         <= #TCQ 1'b0;
      single_cycle_stg2        <= #TCQ 1'b0;
      first_beat_stg2          <= #TCQ 1'b1;
      lower_padded_stg2        <= #TCQ 1'b0;
      lower_padded_stg2_spec   <= #TCQ 1'b0;
      pr_detect_stg2           <= #TCQ 1'b0;
      pr_detect_lanes_stg2     <= #TCQ 2'h0;
      pna_detect_stg2          <= #TCQ 1'b0;
      lresp_detect_stg2        <= #TCQ 1'b0;
      lreq_in_stat_detect_stg2_bit0 <= #TCQ 1'b0; // new signal RC fix
      lreq_in_stat_detect_stg2_bit1 <= #TCQ 1'b0; // new signal RC fix
    end else begin
      // from previous stag_spec
      PR_rcvd_pa_or_pna        <= #TCQ (|pa_detect_stg1 || |pna_detect_stg1) && !prx_in_recoverable_detect;
      data_vld_stg2            <= #TCQ qualified_data_vld_stg1 ||
                                       (data_vld_stg2 && !framing_end_stg2) && rt_stream_enable_stg2;
      in_packet_stg2           <= #TCQ |in_packet_stg1;
      framing_start_stg2       <= #TCQ framing_start_stg1;
      framing_end_stg2         <= #TCQ framing_end_stg1;
      framing_dsc_stg2         <= #TCQ framing_dsc_stg1 || |prx_cs_crc_check_fail[3:2] ||
                                       (prx_cs_crc_check_fail[1] && pd_flag_stg1[0]) || prx_cs_crc_check_fail[0];
      framing_dsc_stg3         <= #TCQ framing_dsc_stg2; // delay framing_dsc, RC fix
      cause_stg2               <= #TCQ cause_stg1;
      //lreq_in_stat_detect_stg2 <= #TCQ !prx_cs_crc_check_fail[2] && !prx_cs_in_error_cond && // org logic
      lreq_in_stat_detect_stg2 <= #TCQ !prx_cs_crc_check_fail[2]
                                       &&
                                       !((prx_cs_in_error_cond  && !PRD_idle2_selected && input_error_state)
                                         && !((|eop_q && ~|  in_packet_stg1))
                                         )
                                         &&     // fix for CR 824086
                                       ((lreq_in_stat_detect_stg1[0] && !prx_cs_crc_check_fail[1]) ||
                                        (lreq_in_stat_detect_stg1[1] && !prx_cs_crc_check_fail[0]))
                                       && // CR# 826090 updates
                                       !(
                                                         PRD_idle2_selected
                                                             &&
                                                         (control_sym_in_error_cond_cmb || idle2_7_4_beat_err_cmb)
                                                            )// CR# 826090 updates, added idle2_7_4_beat_err_cmb in OR condition to fix CR# 849824
                                        ;
      lreq_in_stat_detect_stg2_bit0 <= #TCQ !prx_cs_crc_check_fail[2] && !((prx_cs_in_error_cond  && !PRD_idle2_selected && input_error_state) && !((|eop_q && ~|  in_packet_stg1))) &&   // fix for CR 824086
                                       (lreq_in_stat_detect_stg1[0] && !prx_cs_crc_check_fail[1]); // new logic RC fix

      lreq_in_stat_detect_stg2_bit1 <= #TCQ !prx_cs_crc_check_fail[2] && !((prx_cs_in_error_cond  && !PRD_idle2_selected && input_error_state) && !((|eop_q && ~|  in_packet_stg1))) &&   // fix for CR 824086
                                        (lreq_in_stat_detect_stg1[1] && !prx_cs_crc_check_fail[0]); // new logic RC fix

      PR_phy_rcvd_buf_stat[5]  <= #TCQ (!prx_cs_crc_check_fail[3] && !prx_cs_in_error_cond) ?
                                        (PRD_idle2_selected ? buf_status_stg2[5] : &buf_status_stg2[4:0]) :
                                        PR_phy_rcvd_buf_stat[5];
      PR_phy_rcvd_buf_stat[4:0] <= #TCQ (!prx_cs_crc_check_fail[3] && !prx_cs_in_error_cond) ? buf_status_stg2[4:0] :
                                                                                           PR_phy_rcvd_buf_stat[4:0];
      // from data formatter
      user_def_stg2            <= #TCQ user_def_stg1;
      carryover_stg2           <= #TCQ carryover_stg1;
      // mid_crc_loc_stg2         <= #TCQ mid_crc_loc_stg1; // org logic
      mid_crc_loc_stg2         <= #TCQ mid_crc_loc_stg1 && !PR_phyr_tlast;  // 09_29(2) new logic RC fix
      single_cycle_stg2        <= #TCQ single_cycle_stg1;
      first_beat_stg2          <= #TCQ first_beat_stg1;
      lower_padded_stg2_spec   <= #TCQ lower_padded_stg1 && !framing_end_stg1;
      lower_padded_stg2        <= #TCQ (lower_padded_stg1 && framing_end_stg1) || lower_padded_stg2_spec;
      pr_detect_stg2           <= #TCQ pr_detect_stg1 && ~|prx_cs_crc_check_fail[2:0];
      pr_detect_lanes_stg2     <= #TCQ {2{!prx_cs_crc_check_fail[2]}} &
                                       {(pr_detect_lanes_stg1[1] && !prx_cs_crc_check_fail[0]),
                                        (pr_detect_lanes_stg1[0] && !prx_cs_crc_check_fail[1])};
      pna_detect_stg2          <= #TCQ pna_detect_stg1 && ~|prx_cs_crc_check_fail[2:0];
      lresp_detect_stg2        <= #TCQ !prx_cs_crc_check_fail[2] &&
                                       ((lresp_detect_stg1[1] && !prx_cs_crc_check_fail[0]) ||
                                        (lresp_detect_stg1[0] && !prx_cs_crc_check_fail[1]));
    end
  end

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      buf_status_stg2 <= #TCQ 6'h00;
    end else if (update_buf_stat_stg1 && ~|prx_cs_crc_check_fail[2:0] && !prx_cs_in_error_cond) begin
      buf_status_stg2 <= #TCQ buf_status_stg1;
    end else if (prx_cs_crc_check_fail[3]) begin
      buf_status_stg2 <= #TCQ PR_phy_rcvd_buf_stat;
    end
  end

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      crc_loc_stg2             <= #TCQ 4'b0001;
    end else if (mid_crc_loc_stg1 || !beat_count_q_is_10) begin
      crc_loc_stg2             <= #TCQ crc_loc_stg1;
    end
  end

  // Data gets latched only when both the upper and lower are valid.
  // From this point on, push only complete data fields forward.
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      ordered_rx_data_stg2 <= #TCQ 64'b0;
      vc_stg2              <= #TCQ 1'b0;
      crf_stg2             <= #TCQ 1'b0;
    end else if (qualified_data_vld_stg1) begin
      ordered_rx_data_stg2 <= #TCQ ordered_rx_data_stg1;
      vc_stg2              <= #TCQ vc_stg1;
      crf_stg2             <= #TCQ crf_stg1;
    end
  end

  // take the partial EOP generation from the previous stage and
  // add the consideration for the times when EOP must advance by a cycle
  // when eop_delay is asserted, we could actually send tlast a cycle earlier
  // but we have to wait for the crc check to complete
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      set_eop_stg2     <= #TCQ 1'b0;
      eop_delay_stg2   <= #TCQ 1'b0;
      set_dsc_stg2     <= #TCQ 1'b0;
      dsc_delay_stg2   <= #TCQ 1'b0;
    end else if (!carryover_stg1 && qualified_data_vld_stg1 && !data_vld_stg0[1] && framing_end_stg0) begin
      set_eop_stg2     <= #TCQ 1'b0;
      eop_delay_stg2   <= #TCQ data_stream_enable_stg1;
      set_dsc_stg2     <= #TCQ 1'b0;
      dsc_delay_stg2   <= #TCQ framing_dsc_stg0;
    end else begin
      set_eop_stg2     <= #TCQ (eop_partial_stg1 || eop_delay_stg2) && data_stream_enable_stg1;
      eop_delay_stg2   <= #TCQ 1'b0;
      set_dsc_stg2     <= #TCQ dsc_partial_stg1 || dsc_delay_stg2;
      dsc_delay_stg2   <= #TCQ 1'b0;
    end
  end


  // Generate the destination discontinue signal -
  assign dest_dsc_stg2 = !BR_phyr_tready && PR_phyr_tvalid && data_vld_stg2 &&
                         (!(crc_loc_stg2 == 4'h8) &&
                          !(crc_loc_stg2 == 4'h4 && (mid_crc_loc_stg1 || large_packet_stg3)));


  // }}} End of Stage2 Pipeline Registers -


  // {{{ + Output Error and Retry Handler ---
  reg   [5:0]  output_error_cs;         // Current state of the Output Error Handler
  reg   [5:0]  output_error_ns;         // Next state of the Output Error Handler
  reg          pr_phy_rewind_d;         // Combinatorial rewind
  reg          short_rewind_pulse_d;    // Signal to make rewind assert for only 2 cycles on retry
  reg          short_rewind_pulse;      // Signal to make rewind assert for only 2 cycles on retry
  reg          pr_send_lreq_d;          // Combinatorial Send Link-Request
  reg          pr_send_rfr_d;           // Combinatorial Send Restart-From-Retry
  reg          pr_output_retry_stop_d;  // Indicator that OLLM RX is currently in Output Retry Stopped State
  reg          pr_output_error_stop_d;  // Indicator that OLLM RX is currently in Output Error Stopped State
  reg          pr_port_error_d;         // Indicator that OLLM RX is currently in Port Error State

  // Output Error FSM -
  // Interpretation and combination of the Output error and retry FSMs
  // in Appendix C of the SRIO PHY specification
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      output_error_cs <= #TCQ OUT_RECOVERY_DISABLED;
    end else if (!PR_link_initialized) begin
      output_error_cs <= #TCQ OUT_RECOVERY_DISABLED;
    end else begin
      output_error_cs <= #TCQ output_error_ns;
    end
  end

//--------------------------------------------------------------------------------
  `ifdef SIMULATION

    reg [25*8-1:0] op_err_handler_cs_string = "INVALID";
    reg [25*8-1:0] op_err_handler_ns_string = "INVALID";

    always @* begin
      //output_error_cs
      case (output_error_cs)
        OUT_RECOVERY_DISABLED : op_err_handler_cs_string = "OUT_RECOVERY_DISABLED";
            OUT_WAIT_FOR_EVENT    : op_err_handler_cs_string = "OUT_WAIT_FOR_EVENT";
            OUT_STOP_ERROR        : op_err_handler_cs_string = "OUT_STOP_ERROR";
            OUT_ERROR_RECOVER     : op_err_handler_cs_string = "OUT_ERROR_RECOVER";
            OUT_STOP_RETRY        : op_err_handler_cs_string = "OUT_STOP_RETRY";
            OUT_FATAL             : op_err_handler_cs_string = "OUT_FATAL";
        default               : op_err_handler_cs_string = "INVALID";
      endcase

      //output_error_ns
      case (output_error_ns)
        OUT_RECOVERY_DISABLED : op_err_handler_ns_string = "OUT_RECOVERY_DISABLED";
            OUT_WAIT_FOR_EVENT    : op_err_handler_ns_string = "OUT_WAIT_FOR_EVENT";
            OUT_STOP_ERROR        : op_err_handler_ns_string = "OUT_STOP_ERROR";
            OUT_ERROR_RECOVER     : op_err_handler_ns_string = "OUT_ERROR_RECOVER";
            OUT_STOP_RETRY        : op_err_handler_ns_string = "OUT_STOP_RETRY";
            OUT_FATAL             : op_err_handler_ns_string = "OUT_FATAL";
        default               : op_err_handler_ns_string = "INVALID";
      endcase
     end
  `endif
//--------------------------------------------------------------------------------

  always @* begin
    output_error_ns        = output_error_cs;
    pr_phy_rewind_d        = 1'b0;
    pr_send_lreq_d         = 1'b0;
    pr_send_rfr_d          = 1'b0;
    short_rewind_pulse_d   = 1'b0;
    pr_output_retry_stop_d = 1'b0;
    pr_output_error_stop_d = 1'b0;
    pr_port_error_d        = 1'b0;

    case (output_error_cs)
    OUT_RECOVERY_DISABLED : begin
      if (PR_link_initialized) begin
        output_error_ns        = OUT_WAIT_FOR_EVENT;
      end
    end

    OUT_WAIT_FOR_EVENT : begin
      if (prx_out_fatal_detect) begin
        output_error_ns        = OUT_FATAL;
        pr_phy_rewind_d        = 1'b1;
      end else if ((pna_detect_stg2 && !prx_cs_crc_check_fail[3]) || prx_out_recoverable_detect) begin
        output_error_ns        = OUT_STOP_ERROR;
        pr_phy_rewind_d        = 1'b1;
      end else if (pr_detect_stg2 && !prx_cs_crc_check_fail[3]) begin
        output_error_ns        = OUT_STOP_RETRY;
        short_rewind_pulse_d   = 1'b1; // makes rewind only assert for 2 cycles on a retry event
        pr_phy_rewind_d        = 1'b1;
      end
    end

    OUT_STOP_ERROR : begin
      pr_phy_rewind_d        = 1'b1;
      pr_send_lreq_d         = 1'b1;
      pr_output_error_stop_d = 1'b1;
      if (prx_out_fatal_detect) begin
        output_error_ns        = OUT_FATAL;
        pr_send_lreq_d         = 1'b0;
      end else if (PT_lreq_sent) begin
        output_error_ns        = OUT_ERROR_RECOVER;
        pr_send_lreq_d         = 1'b0;
      end
    end

    OUT_ERROR_RECOVER: begin
      pr_phy_rewind_d        = 1'b1;
      pr_output_error_stop_d = 1'b1;
      if (prx_out_fatal_detect) begin
        output_error_ns        = OUT_FATAL;
      end else if (lresp_detect_stg3 && ((|pr_detect_lanes_stg3[0]) ||
                                         (pr_detect_stg2 && !prx_cs_crc_check_fail[3]))) begin
        output_error_ns        = OUT_STOP_RETRY;
        short_rewind_pulse_d   = 1'b1; // makes rewind only assert for 2 cycles on a retry event
        pr_phy_rewind_d        = 1'b1;
      end else if (prx_force_send_lreq) begin
        output_error_ns        = OUT_STOP_ERROR;
      end else if (lresp_detect_stg3) begin
        output_error_ns        = OUT_WAIT_FOR_EVENT;
      end
    end

    OUT_STOP_RETRY : begin
      pr_send_rfr_d          = !(pna_detect_stg1 || prx_out_recoverable_detect);
      pr_send_lreq_d         = (pna_detect_stg1 || prx_out_recoverable_detect);
      pr_phy_rewind_d        = short_rewind_pulse;
      pr_output_retry_stop_d = !(pna_detect_stg1 || prx_out_recoverable_detect);
      pr_output_error_stop_d = (pna_detect_stg1 || prx_out_recoverable_detect);
      if (prx_out_fatal_detect) begin
        output_error_ns        = OUT_FATAL;
      end else if (pna_detect_stg1 || prx_out_recoverable_detect) begin
        pr_phy_rewind_d        = 1'b1;
        output_error_ns        = OUT_STOP_ERROR;
      end else if (PT_rfr_sent) begin
        output_error_ns        = OUT_WAIT_FOR_EVENT;
        pr_send_rfr_d          = 1'b0;
      end
    end

    OUT_FATAL : begin
      pr_phy_rewind_d        = 1'b1;
      pr_port_error_d        = 1'b1;
      if (PC_clr_port_error) begin
        output_error_ns        = OUT_RECOVERY_DISABLED;
      end
    end

    default : begin
      output_error_ns        = OUT_FATAL;
      pr_phy_rewind_d        = 1'b1;
      pr_port_error_d        = 1'b1;
    end
    endcase
  end

  // Drive output control signals to OLLM TX
  reg pc_load_ackids_q;
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PR_rewind            <= #TCQ 1'b0;
      PR_send_lreq         <= #TCQ 1'b0;
      PR_send_rfr          <= #TCQ 1'b0;
      PR_output_retry_stop <= #TCQ 1'b0;
      PR_output_error_stop <= #TCQ 1'b0;
      PR_port_error        <= #TCQ 1'b0;
      short_rewind_pulse   <= #TCQ 1'b0;
      pc_load_ackids_q     <= #TCQ 1'b0;
    end else begin
      PR_rewind            <= #TCQ pr_phy_rewind_d || (PC_load_ackids || pc_load_ackids_q);
      PR_send_lreq         <= #TCQ pr_send_lreq_d;
      PR_send_rfr          <= #TCQ pr_send_rfr_d;
      PR_output_retry_stop <= #TCQ pr_output_retry_stop_d;
      PR_output_error_stop <= #TCQ pr_output_error_stop_d;
      PR_port_error        <= #TCQ pr_port_error_d;
      short_rewind_pulse   <= #TCQ short_rewind_pulse_d;
      pc_load_ackids_q     <= #TCQ PC_load_ackids;
    end
  end


    // *- COVERAGE (cp_PR_pr_and_pna_same_cycle)
    // Observe pr_detect_stg1 and pna_detect_stg1 on the same cycle

    // *- COVERAGE (cp_PR_pr_1before_pna)
    // Observe pr_detect_stg1 one cycle before pna_detect_stg1

    // *- COVERAGE (cp_PR_pr_2before_pna)
    // Observe pr_detect_stg1 two cycles before pna_detect_stg1

    // *- COVERAGE (cp_PR_pr_3before_pna)
    // Observe pr_detect_stg1 three cycles before pna_detect_stg1

    // *- COVERAGE (cp_PR_pna_1before_pr)
    // Observe pna_detect_stg1 one cycle before pr_detect_stg1

    // *- COVERAGE (cp_PR_pna_2before_pr)
    // Observe pna_detect_stg1 two cycles before pr_detect_stg1

    // *- COVERAGE (cp_PR_pna_3before_pr)
    // Observe pna_detect_stg1 three cycles before pr_detect_stg1

    // *- COVERAGE (cp_PR_link_init_cross_output_fsm)
    // Observe link_initialized deassert while the Output Error and
    // Retry fsm is in each and every state


  // }}} end of Output Error and Retry ----


  // {{{ + Input Error and Retry Handler ----
  reg   [6:0]  input_error_cs;          // Current state of the Input Error Handler
  reg   [6:0]  input_error_ns;          // Next state of the Input Error Handler
  reg          pr_send_pna_early;       // Combinatorial Send Packet-Not_Accepted - early
  reg          pr_send_pna_early_q;     // Combinatorial Send Packet-Not_Accepted - early reg
  reg          pr_send_pna_d;           // Combinatorial Send Packet-Not_Accepted
  reg          pr_send_pr_early;        // Combinatorial Send Packet-Retry - early
  reg          pr_send_pr_early_q;      // Combinatorial Send Packet-Retry - early reg
  reg          pr_send_pr_d;            // Combinatorial Send Packet-Retry
  reg          pr_send_lresp_d;         // Combinatorial Send Link-Response
  reg          pr_input_retry_stop_d;   // Indicator that OLLM RX is currently in Input Retry Stopped State
  reg          pr_input_error_stop_d;   // Indicator that OLLM RX is currently in Input Error Stopped State
  reg          pr_input_status_good_d;  // Indicator that OLLM RX is currently in Input Waiting for Event State
  reg   [4:0]  pr_port_stat_early;      // Current port status
  reg   [4:0]  pr_port_stat_early_q;    // Current port status
  reg   [4:0]  pr_port_stat_d;          // Current port status
  reg          rt_stream_enable_stg2_d; // Combinatorial, Used to enable the stream for RT
  reg          mask_crc_error_d;        // mask an error on the same beat as a lresp
  reg          mask_crc_error;          // mask an error on the same beat as a lresp
  reg   [3:0]  prx_cs_crc_check_fail_q; // used to generate cs_crc_in_error_cond
  reg          delayed_error_detect_d;  // used when there is an error detected between LREQ (rcvd) and LRESP (sent)
  reg          delayed_error_detect;    // used when there is an error detected between LREQ (rcvd) and LRESP (sent)
  reg          set_port_stat_ok;        // added to fix CR# 822469
  reg          set_port_stat_ok_q;      // added to fix CR# 822469
  reg          multi_lreq;              // new signal declaration RC fix
  reg          multi_lreq_q;                // new signal RC fix
  reg          lreq_recov_err;          // new signal RC fix
  reg          lreq_recov_err_q;        // new signal RC fix

//---------- Display the input error port recovery and retry states ----
  `ifdef SIMULATION  // While fixing CR# 822469, added below display comments for easy debug

    reg [25*8-1:0] ip_err_handler_cs_string = "INVALID";
    reg [25*8-1:0] ip_err_handler_ns_string = "INVALID";

    always @* begin
    //input_error_cs
    case (input_error_cs)
    IN_RECOVERY_DISABLED  : ip_err_handler_cs_string = "IN_RECOVERY_DISABLED";
        IN_WAIT_FOR_EVENT     : ip_err_handler_cs_string = "IN_WAIT_FOR_EVENT";
        IN_STOP_INPUT         : ip_err_handler_cs_string = "IN_STOP_INPUT";
        IN_ERROR_STOPPED      : ip_err_handler_cs_string = "IN_ERROR_STOPPED";
        IN_ERROR_RECOVERY     : ip_err_handler_cs_string = "IN_ERROR_RECOVERY";
        IN_RETRY_STOPPED      : ip_err_handler_cs_string = "IN_RETRY_STOPPED";
        IN_REC_DISABLED_LRESP : ip_err_handler_cs_string = "IN_REC_DISABLED_LRESP";
    default               : ip_err_handler_cs_string = "INVALID";
    endcase

    //input_error_ns
    case (input_error_ns)
    IN_RECOVERY_DISABLED  : ip_err_handler_ns_string = "IN_RECOVERY_DISABLED";
        IN_WAIT_FOR_EVENT     : ip_err_handler_ns_string = "IN_WAIT_FOR_EVENT";
        IN_STOP_INPUT         : ip_err_handler_ns_string = "IN_STOP_INPUT";
        IN_ERROR_STOPPED      : ip_err_handler_ns_string = "IN_ERROR_STOPPED";
        IN_ERROR_RECOVERY     : ip_err_handler_ns_string = "IN_ERROR_RECOVERY";
        IN_RETRY_STOPPED      : ip_err_handler_ns_string = "IN_RETRY_STOPPED";
        IN_REC_DISABLED_LRESP : ip_err_handler_ns_string = "IN_REC_DISABLED_LRESP";
    default               : ip_err_handler_ns_string = "INVALID";
    endcase

    end
  `endif
//--------------------------------------------------------------------------------
  `ifdef SIMULATION

    reg [25*8-1:0] pr_port_stat_string = "PORT_STAT_OK";

    always @* begin
      //output_error_cs
      case (pr_port_stat_d)
        PORT_STAT_ERROR      : pr_port_stat_string = "PORT_STAT_ERROR     ";
        PORT_STAT_RETRY_STOP : pr_port_stat_string = "PORT_STAT_RETRY_STOP";
        PORT_STAT_ERROR_STOP : pr_port_stat_string = "PORT_STAT_ERROR_STOP";
        PORT_STAT_OK         : pr_port_stat_string = "PORT_STAT_OK        ";
        default              : pr_port_stat_string = "PORT_STAT_OK        ";
      endcase
     end
  `endif
//--------------------------------------------------------------------------------

  // Input Error FSM -
  // Interpretation and combination of the Input error and retry FSMs
  // in Appendix C of the SRIO PHY specification
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      input_error_cs <= #TCQ IN_RECOVERY_DISABLED;
    end else if (!PP_port_initialized) begin
      input_error_cs <= #TCQ IN_RECOVERY_DISABLED;
    end else begin
      input_error_cs <= #TCQ input_error_ns;
    end
  end

  // when core is in error recovery state and SOP + LREQ comes in b2b packets, then detect
  // LREQ. so use below signal to make the lreq_in_stat_detect_stg2 active
  // (as lreq_in_stat_detect_stg1 would have been active)
  assign input_error_state = (input_error_cs == IN_ERROR_STOPPED) ? 1'b0 : 1'b1;

  // when core is in error recovery state and SOP + LREQ comes in b2b packets, then detect
  // LREQ. so use below signal to make the lreq_in_stat_detect_stg2 active
  // (as lreq_in_stat_detect_stg1 would have been active)
  assign in_retry_stopped_state = (input_error_cs == IN_RETRY_STOPPED) ? 1'b1 : 1'b0;
  assign not_in_retry_stopped_state = (input_error_ns == IN_RETRY_STOPPED) ? 1'b0 : 1'b1;

  // added below condition to fix the CR# 837481 //
  assign in_error_stopped_state = (input_error_cs == IN_ERROR_STOPPED) ? 1'b1 : 1'b0;

reg no_lresp_sending;
reg no_lresp_sending_stg0;

  always @* begin
    input_error_ns          = input_error_cs;
    pr_send_pna_early       = 1'b0;
    pr_send_pna_d           = 1'b0;
    pr_send_pr_early        = 1'b0;
    pr_send_pr_d            = 1'b0;
    pr_send_lresp_d         = 1'b0;
    rt_stream_enable_stg2_d = 1'b0;
    pr_input_retry_stop_d   = 1'b0;
    pr_input_error_stop_d   = 1'b0;
    pr_input_status_good_d  = 1'b0;
    delayed_error_detect_d  = 1'b0;
    mask_crc_error_d        = 1'b0;
    set_port_stat_ok        = 1'b0;// added as switch to fix CR# 822469
    multi_lreq              = 1'b0;// default assignment, new logic, RC fix
    lreq_recov_err          = 1'b0;// default assignment, new logic, RC fix
    pr_port_stat_d          = PORT_STAT_OK;
    pr_port_stat_early      = PORT_STAT_OK;
    no_lresp_sending        = 1'b0;

    case (input_error_cs)
    IN_RECOVERY_DISABLED : begin
      rt_stream_enable_stg2_d  = PR_link_initialized && PC_error_disable;
      // still must respond to a LREQ, even if FSM is disabled
      if (lreq_in_stat_detect_stg2 && !prx_cs_crc_check_fail[3]) begin
        input_error_ns          = IN_REC_DISABLED_LRESP;
      end else if (PR_link_initialized && !PC_error_disable) begin
        input_error_ns          = IN_WAIT_FOR_EVENT;
      end
    end

    IN_WAIT_FOR_EVENT : begin
      rt_stream_enable_stg2_d = 1'b1;
      pr_input_status_good_d  = 1'b1;
      //if (enable_state_stg1 && (prx_in_recoverable_detect || prx_in_retry_detect)) begin // fix for 821477
      //if (enable_state_stg1 && (prx_in_recoverable_detect || prx_in_retry_detect) && !lreq_in_stat_detect_stg2) begin // fix for 821477 updated logic
      if (enable_state_stg1 && (prx_in_recoverable_detect || prx_in_retry_detect) && !lreq_in_stat_detect_stg2_bit0) begin // fix for 821477, new fix for few issues, RC fix
          input_error_ns          = IN_STOP_INPUT;
          rt_stream_enable_stg2_d = 1'b0;
          pr_send_pna_early       = prx_in_recoverable_detect || !RETRY;
          pr_send_pr_early        = prx_in_retry_detect && !prx_in_recoverable_detect && RETRY;
              if (lreq_in_stat_detect_stg2_bit1 && !prx_cs_crc_check_fail[3]) begin
                  lreq_recov_err = 1'b1;// to detect lreq, new logic
              end
      end else if (lreq_in_stat_detect_stg2 && !prx_cs_crc_check_fail[3]) begin
        // added set_port_stat_ok as switch (or flag) here to fix CR# 822469
        // When in WAIT_FOR_EVENT state, if recoverable error occurs, then pass this error bit as port status
            set_port_stat_ok        = prx_in_recoverable_detect;// added to fix CR# 822469
        input_error_ns          = IN_ERROR_RECOVERY;
      end
    end

    IN_STOP_INPUT : begin
      pr_send_pna_d           = pr_send_pna_early_q || PR_send_pna || prx_in_recoverable_detect;
      pr_send_pr_d            = ((pr_send_pr_early_q && !prx_in_recoverable_detect) || PR_send_pr) && !PT_pr_sent;
      pr_port_stat_d          = pr_send_pna_d ? PORT_STAT_ERROR_STOP : PORT_STAT_RETRY_STOP;
   //   multi_lreq              = multi_lreq_q;
      lreq_recov_err          = lreq_recov_err_q; // new logic to keep the lreq_recov_err registered value
      //if ((lreq_in_stat_detect_stg2 && !prx_cs_crc_check_fail[3]) || delayed_error_detect) begin // org logic
      if ((lreq_in_stat_detect_stg2 && !prx_cs_crc_check_fail[3]) || delayed_error_detect || lreq_recov_err) begin // updated to fix the delayed_error_detect.
        delayed_error_detect_d  = 1'b1;
      end
      // this is the case where we are in retry but we receive a LREQ
      //if ((PT_pr_sent || PT_pna_sent) && // org logic
          //(delayed_error_detect || (lreq_in_stat_detect_stg2 && !prx_cs_crc_check_fail[3]))) begin // org logic
      if (((PT_pr_sent || PT_pna_sent) && // new logic
          (delayed_error_detect || (lreq_in_stat_detect_stg2 && !prx_cs_crc_check_fail[3]))) || multi_lreq) begin   // 09_30(2) new logic
        input_error_ns          = IN_ERROR_RECOVERY;
        mask_crc_error_d        = |prx_cs_crc_check_fail_q[2:0];
        rt_stream_enable_stg2_d = 1'b1;
        delayed_error_detect_d  = 1'b0;
        pr_send_pna_d           = 1'b0;
        pr_send_pr_d            = 1'b0;
        pr_port_stat_early      = pr_port_stat_d; // PR_port_stat;//
        lreq_recov_err          = 1'b0; // force the lre_recovery error to 0, newly added
        //no_lresp_sending        = 1'b1;
      end else if (PT_pna_sent) begin
        input_error_ns          = IN_ERROR_STOPPED;
        pr_send_pna_d           = 1'b0;
        pr_send_pr_d            = 1'b0;
      end else if (!pr_send_pna_d && PT_pr_sent && RETRY) begin
        input_error_ns          = IN_RETRY_STOPPED;
        pr_send_pr_d            = 1'b0;
      end
    end

    IN_ERROR_STOPPED : begin
      pr_input_error_stop_d   = 1'b1;
      pr_port_stat_d          = PORT_STAT_ERROR_STOP;
      pr_port_stat_early      = PORT_STAT_ERROR_STOP;

   // commented below logic as from ERROR STOPPED state, only way to get out is in ERROR RECOVERY state.
   //   if (lreq_in_stat_detect_stg2 && !prx_cs_crc_check_fail[3] &&
   //       (prx_in_recoverable_detect || prx_in_retry_detect) && !pp_out_of_sync_stg1) begin
   //     pr_send_pna_early       = prx_in_recoverable_detect || pr_send_pna_early_q;
   //     pr_send_pr_early        = prx_in_retry_detect || pr_send_pr_early_q;
   //     rt_stream_enable_stg2_d = 1'b0;
   //     input_error_ns          = IN_STOP_INPUT;
   //   end else if (lreq_in_stat_detect_stg2 && !prx_cs_crc_check_fail[3]) begin
      if (lreq_in_stat_detect_stg2 && !prx_cs_crc_check_fail[3]) begin
        input_error_ns          = IN_ERROR_RECOVERY;
        mask_crc_error_d        = |prx_cs_crc_check_fail_q[2:0];
        rt_stream_enable_stg2_d = 1'b1;
            if (prx_in_recoverable_detect && lreq_in_stat_detect_stg2_bit1) begin // newly added
                lreq_recov_err = 1'b1;
            end
      end
    end

    IN_ERROR_RECOVERY : begin
      pr_input_error_stop_d   = 1'b0;
//    pr_send_lresp_d         = !in_packet_stg3;// deactivated signal behavior
      rt_stream_enable_stg2_d = 1'b1;
      pr_input_status_good_d  = 1'b1;
      multi_lreq              = 1'b0;            // new addition
      lreq_recov_err          = lreq_recov_err_q;// new addition
      set_port_stat_ok        = set_port_stat_ok_q;     //

      if (!PR_phyr_tvalid && !PR_phyr_tlast && !pr_phyr_tlast_d) begin
                                 // if there is no PD error in LREQ, then only generate the LRESP
         pr_send_lresp_d         = !lreq_pd_error;  // CR 825487 logic updates
         // old logic before 27 nov
         //pr_send_lresp_d         = !lreq_pd_error;//1'b1;              // 09_30(3), newly added
      end else begin
         pr_send_lresp_d         = PR_send_lresp;      // 09_30(3), newly added
      end

      //if (set_port_stat_ok || idle_seq_in_error_cond_cmb) begin                       // added as switch to fix CR# 822469
      if (set_port_stat_ok) begin                       // added as switch to fix CR# 822469
        pr_port_stat_d          = PORT_STAT_ERROR_STOP; // If the state machine is coming from IN_WAIT_FOR_EVENT state
        pr_port_stat_early      = PORT_STAT_ERROR_STOP; // and if the recoverable error occurs in that state, then
      end else begin                                                    // generate port status as ERROR STOPPED
        pr_port_stat_d          = pr_port_stat_early_q; // else pass the present state of the port status
        pr_port_stat_early      = pr_port_stat_early_q; // as is.
      end                                                                       //
 //     if ((lreq_in_stat_detect_stg2 && !prx_cs_crc_check_fail[3]) || prx_in_retry_detect || delayed_error_detect) begin   // 09_30(2) org logic
 //     if ((prx_in_recoverable_detect && !mask_crc_error) || prx_in_retry_detect || delayed_error_detect) begin // updated logic
      if ((prx_in_recoverable_detect && !mask_crc_error && !prx_in_recoverable_detect_delay)
          ||                                             // CR# 851432 fixed by adding !prx_in_recoverable_detect_delay in above statement
          prx_in_retry_detect
          ||
          delayed_error_detect
          ||
          lreq_recov_err) begin
        delayed_error_detect_d  = !PT_lresp_sent
                                  &&              // Added to fix the CR 825487
                                  !lreq_pd_error; // when LREQ PD error present, dont detect any
                                                  // other error when core is in IN_ERROR_RECOVERY state
                                                  // wait for clear LREQ.
        pr_send_pna_early       = prx_in_recoverable_detect || pr_send_pna_early_q || lreq_recov_err; // updated PNA sending logic
        pr_send_pr_early        = prx_in_retry_detect || pr_send_pr_early_q;                          // updated PR sending logic
 //     pr_send_pna_early       = prx_in_recoverable_detect || pr_send_pna_early_q;
 //     pr_send_pr_early        = prx_in_retry_detect || pr_send_pr_early_q;
 //     pr_send_pna_early       = 1'b0;  // fix for CR 797396, negated pna sending
 //     pr_send_pr_early        = 1'b0;
          lreq_recov_err        = 1'b0;// disabled the lreq recovery error
      end
   //   if (( prx_in_retry_detect || delayed_error_detect) &&                          // 09_30(2)
      if (((prx_in_recoverable_detect && !mask_crc_error) || prx_in_retry_detect || delayed_error_detect) &&   // 09_30(2)
        enable_state_stg1 && PT_lresp_sent) begin
        pr_send_pna_early       = prx_in_recoverable_detect || pr_send_pna_early_q;
        pr_send_pr_early        = prx_in_retry_detect || pr_send_pr_early_q;
        rt_stream_enable_stg2_d = 1'b0;
        pr_send_lresp_d         = 1'b0;
        set_port_stat_ok        = 1'b0; // reset the switch while exiting this state, added to fix CR# 822469
//      multi_lreq              = 1'b1;
        input_error_ns          = IN_STOP_INPUT;
        //no_lresp_sending        = 1'b0;
      end else if (PT_lresp_sent) begin
        pr_send_lresp_d         = 1'b0;
        set_port_stat_ok            = 1'b0; // reset the switch while exiting this state, added to fix CR# 822469
        input_error_ns          = IN_WAIT_FOR_EVENT;
        //no_lresp_sending        = 1'b0;
      end
    end

    IN_REC_DISABLED_LRESP : begin // only hit when LREQ is received when FSM is disabled
      pr_send_lresp_d         = 1'b1;
      if (PT_lresp_sent) begin
        pr_send_lresp_d         = 1'b0;
        input_error_ns          = IN_RECOVERY_DISABLED;
      end
    end

    IN_RETRY_STOPPED : begin
      pr_port_stat_d          = PORT_STAT_RETRY_STOP;
      pr_input_retry_stop_d   = 1'b1;
      rt_stream_enable_stg2_d = |rfr;
      // always need to be able to detect an error, even when servicing a retry
      if (enable_state_stg1) begin
        if (prx_in_recoverable_detect) begin
          pr_send_pna_early       = 1'b1;
          input_error_ns          = IN_STOP_INPUT;
        end else if (lreq_in_stat_detect_stg2 && !prx_cs_crc_check_fail[3]) begin
          input_error_ns          = IN_ERROR_RECOVERY;
          mask_crc_error_d        = |prx_cs_crc_check_fail_q[2:0];
          rt_stream_enable_stg2_d = 1'b1;
          pr_port_stat_early      = PORT_STAT_RETRY_STOP;// Added to send the port status as 5
                                                         // while entering in the error recovery state
        end else if (rfr_detect_stg1) begin
          input_error_ns          = IN_WAIT_FOR_EVENT;
          pr_port_stat_d          = PORT_STAT_OK;
          pr_input_status_good_d  = 1'b1;
          rt_stream_enable_stg2_d = 1'b1;
        end
      end
    end

    default : begin
      input_error_ns          = IN_RECOVERY_DISABLED;
    end
    endcase
  end

  // Drive input control signals to OLLM TX
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      pr_send_pna_early_q     <= #TCQ 1'b0;
      PR_send_pna             <= #TCQ 1'b0;
      pr_send_pr_early_q      <= #TCQ 1'b0;
      PR_send_pr              <= #TCQ 1'b0;
      PR_send_lresp           <= #TCQ 1'b0;
      PR_input_error_stop     <= #TCQ 1'b0;
      PR_input_retry_stop     <= #TCQ 1'b0;
      PR_port_stat            <= #TCQ PORT_STAT_OK;
      pr_port_stat_early_q    <= #TCQ PORT_STAT_OK;
      PR_port_stat_ok         <= #TCQ 1'b1;
      PR_input_status_good    <= #TCQ 1'b0;
      rt_stream_enable_stg2   <= #TCQ 1'b0;
      prx_cs_crc_check_fail_q <= #TCQ 4'h0;
      mask_crc_error          <= #TCQ 1'b0;
      delayed_error_detect    <= #TCQ 1'b0;
      set_port_stat_ok_q      <= #TCQ 1'b0;             // registered version of the switch, added to fix CR# 822469
      multi_lreq_q            <= #TCQ 1'b0;// default values
      err_recovery            <= #TCQ 1'b0;// default values
      lreq_recov_err_q        <= #TCQ 1'b0;// default values
      no_lresp_sending_stg0   <= #TCQ 1'b0;


    end else begin
      pr_send_pna_early_q     <= #TCQ pr_send_pna_early;
      PR_send_pna             <= #TCQ pr_send_pna_d;
      pr_send_pr_early_q      <= #TCQ pr_send_pr_early;
      PR_send_pr              <= #TCQ pr_send_pr_d;
      PR_send_lresp           <= #TCQ pr_send_lresp_d && !PT_lresp_sent;
      PR_input_error_stop     <= #TCQ pr_input_error_stop_d;
      PR_input_retry_stop     <= #TCQ pr_input_retry_stop_d;
      PR_port_stat            <= #TCQ pr_port_stat_d;
      pr_port_stat_early_q    <= #TCQ pr_port_stat_early;
      PR_port_stat_ok         <= #TCQ pr_port_stat_d == PORT_STAT_OK;
      PR_input_status_good    <= #TCQ pr_input_status_good_d;
      rt_stream_enable_stg2   <= #TCQ rt_stream_enable_stg2_d;
      prx_cs_crc_check_fail_q <= #TCQ prx_cs_crc_check_fail;
      mask_crc_error          <= #TCQ mask_crc_error_d;
      delayed_error_detect    <= #TCQ delayed_error_detect_d;
      set_port_stat_ok_q      <= #TCQ set_port_stat_ok;// registered version of the switch, added to fix CR# 822469
      multi_lreq_q            <= #TCQ multi_lreq;      // create one level pipeline
      lreq_recov_err_q        <= #TCQ lreq_recov_err;  // create one level pipeline
      err_recovery            <= #TCQ input_error_ns == IN_ERROR_RECOVERY; // create one level pipeline
      no_lresp_sending_stg0   <= #TCQ no_lresp_sending;
    end
  end


    // *- COVERAGE (cp_PR_error_cross_input_fsm)
    // Observe in_recoverable_detect (input error) assert while the Input Error
    // and Retry fsm is in each of the states

    // *- COVERAGE (cp_PR_rewind_cross_input_fsm)
    // Observe in_retry_detect (input rewind) assert while the Input Error
    // and Retry fsm is in each of the states

    // *- COVERAGE (cp_PR_link_init_cross_input_fsm)
    // Observe PR_link_initialized deassert while the Input Error and Retry
    // fsm is in each and every state

    // *- COVERAGE (cp_PR_error_disable_enumerate)
    // Observe both values of PC_error_disable

    // *- COVERAGE (cp_PR_port_stat_enumerate)
    // Observe the four expected values of PR_port_stat

    // *- ASSERTION (ap_PR_port_status_illegal)
    // PR_port_status will never be Unrecoverable or Reserved

    // *- ASSERTION (ap_PR_send_pna_and_send_pr)
    // PR_send_pna and PR_send_pr should never assert on the same cycle

    // *- COVERAGE (cp_PR_ct_cross_input_fsm)
    // Cross the delivery of continuous traffic packet data with all
    // states of the Input Error state machine

    // *- COVERAGE (cp_PR_stomp_and_stream_enabled)
    // Receive a stomp control symbol while in regular operation

    // *- COVERAGE (cp_PR_stomp_and_stream_disabled)
    // Receive a stomp control symbol while in the stopped state

    // *- COVERAGE (cp_PR_lreq_detected_before_link_initialized)
    // Observe a LREQ when link is not initialized


  // }}} End of Input Error and Retry -----

// }}} End Stage2 Pipeline ---------------


// {{{ Stage3 Pipeline -------------------

  // pipeline registers
  // - This stage constists of a delay stage to allow error detection
  // logic to catch up with the output of the OLLM RX to the Buffer
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      rt_stream_enable_stg3 <= #TCQ 1'b0;
      data_vld_stg3         <= #TCQ 1'b0;
      lresp_detect_stg3     <= #TCQ 1'b0;
      pr_detect_lanes_stg3  <= #TCQ 1'b0;
      //standard_dsc_case_delay  <= #TCQ 1'b0;//CR 821476 removed assignment
      prx_in_recoverable_detect_delay  <= #TCQ 1'b0;//CR 821476
    end else begin
      rt_stream_enable_stg3 <= #TCQ rt_stream_enable_stg2;
      data_vld_stg3         <= #TCQ data_vld_stg2 && (qualified_data_vld_stg1 || framing_end_stg2) &&
                                    !(first_beat_stg2 && framing_dsc_stg2);
      lresp_detect_stg3     <= #TCQ lresp_detect_stg2 && !prx_cs_crc_check_fail[3];
      pr_detect_lanes_stg3  <= #TCQ pr_detect_lanes_stg2 & {2{!prx_cs_crc_check_fail[3]}};
//      standard_dsc_case_delay  <= #TCQ standard_dsc_case;//CR 821476
      prx_in_recoverable_detect_delay  <= #TCQ prx_in_recoverable_detect;//CR 821476
    end
  end

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      in_packet_stg3       <= #TCQ 1'b0;
      ordered_rx_data_stg3 <= #TCQ 64'b0;
      vc_stg3              <= #TCQ 1'b0;
      crf_stg3             <= #TCQ 1'b0;
      dest_dsc_stg3        <= #TCQ 1'b0;
      mid_crc_loc_stg3     <= #TCQ 1'b0;
      set_eop_stg3         <= #TCQ 1'b0;
      set_dsc_stg3         <= #TCQ 1'b0;
      eop_delay_stg3       <= #TCQ 1'b0;
      framing_start_stg3   <= #TCQ 1'b0;
      framing_end_stg3     <= #TCQ 1'b0;
      lower_padded_stg3    <= #TCQ 1'b0;
      single_cycle_stg3    <= #TCQ 1'b0;
    end else if (advance_condition) begin
      in_packet_stg3       <= #TCQ in_packet_stg2;
      ordered_rx_data_stg3 <= #TCQ ordered_rx_data_stg2;
      vc_stg3              <= #TCQ vc_stg2;
      crf_stg3             <= #TCQ crf_stg2;
      dest_dsc_stg3        <= #TCQ dest_dsc_stg2 || framing_dsc_stg2;
      mid_crc_loc_stg3     <= #TCQ mid_crc_loc_stg2;
      set_eop_stg3         <= #TCQ set_eop_stg2;
      set_dsc_stg3         <= #TCQ set_dsc_stg2;
      eop_delay_stg3       <= #TCQ eop_delay_stg2;
      framing_start_stg3   <= #TCQ framing_start_stg2;
      framing_end_stg3     <= #TCQ framing_end_stg2;
      lower_padded_stg3    <= #TCQ lower_padded_stg2;
      single_cycle_stg3    <= #TCQ single_cycle_stg2;
    end
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      crc_loc_stg3         <= #TCQ 4'b0001;
    end else if (advance_condition) begin
      // special case to forward the crc location by one beat for certain types of very small packets
      if (data_vld_stg2 && framing_end_stg2 && framing_start_stg3 && (!data_vld_stg3 || framing_end_stg3)) begin
        crc_loc_stg3         <= #TCQ crc_loc_stg1;
      end else begin
        crc_loc_stg3         <= #TCQ crc_loc_stg2;
      end
    end
  end

  // when asserted, indicates a packet is larger than 80 bytes
  always @(posedge phy_clk) begin
    if (phy_rst_q)
      large_packet_stg3 <= #TCQ 1'b0;
    else if (pr_phyr_tlast_d || PR_input_retry_stop || PR_input_error_stop || PR_send_pna)// added PR_send_pna
      large_packet_stg3 <= #TCQ 1'b0;
  //  else if (mid_crc_loc_stg2 && !mid_crc_loc_stg3) // org logic
    else if ((mid_crc_loc_stg2 && !mid_crc_loc_stg3) && data_vld_stg3)     // 09_30(1) added data valid signal
      large_packet_stg3 <= #TCQ 1'b1;
  end
  // end of pipeline registers

// }}} End Stage3 Pipeline ---------------


// {{{ Stage4 Pipeline -------------------

  // {{{ + RX Buf Interface -----------------
// FIXVC - add VC parameters here
// VC, VC1_CT
  reg       tvalid_delay;
  reg       stalled_discontinue;
  reg       packet_discontinue;
  reg       tlast_on_mid_crc, tlast_on_mid_crc_d;
// NOTE - CFR adding or removing tvalid_delay isn't fixing this. What about observing dsc_partial_stg1 vs
// dsc_delay_stg2? When dsc_delay_stg2 is asserted, 2 cycles before tvalid_delay,
// the equation should be set_dsc_stg3, ignoring tvalid_delay. note that eop_delay_stg2 matches the behavior
// of dsc_delay_stg2.
// When dsc_partial_stg1, ?
  assign      standard_dsc_case = ((dest_dsc_stg3 || set_dsc_stg3) && !(tvalid_delay && !set_eop_stg3))
                                  ||
                                  prx_in_recoverable_detect
                                      // CR 826089, below condition is added to detect the PD errors in
                                  ||  // IDLE2 packets                                 //
                                  (PRD_idle2_selected && control_sym_in_error_cond_cmb)//
                                ;

  assign    advance_condition = BR_phyr_tready || !PR_phyr_tvalid;

  // TLAST generation -
  // Assert TLAST when:
  // 1) CRC is removed and causes the last word to shift by one
  // 2) there is a source or dest discontinue
  // 3) carry forward of partial EOP calculation from stage 2
  // TUSER[0] generation (packet_discontinue) -
  // TUSER is distinct from the other bits, in that it is only driven
  // on TLAST. So, it is driven by the same logic.
  always @* begin
    if (advance_condition) begin
      // don't assert tlast if an error/retry happened before the beginning of a packet
//       if (((out_of_packet && !(PR_phyr_tvalid && BR_phyr_tready)) || // org logic
      if (((out_of_packet && !(PR_phyr_tvalid && BR_phyr_tready)) ||
           (PR_phyr_tvalid && BR_phyr_tready && PR_phyr_tlast)) &&
             (standard_dsc_case || (!vc_stg3 && (!rt_stream_enable_stg3 || !rt_stream_enable_stg2)))) begin
        pr_phyr_tlast_d    = 1'b0;
        tlast_on_mid_crc_d = 1'b0;
        packet_discontinue = 1'b0;
      // last beat is also where the mid-crc should be
      end else if (mid_crc_loc_stg2 && framing_end_stg2 && lower_padded_stg2) begin
        pr_phyr_tlast_d    = 1'b1;
        tlast_on_mid_crc_d = 1'b1;
        packet_discontinue = (standard_dsc_case || framing_dsc_stg2 ||
                              stalled_discontinue || prx_cs_crc_check_fail[3]);
      // early tlast when removing the crc causes a beat to be removed
      end else if (((crc_loc_stg2 == 4'h8) || (crc_loc_stg2 == 4'h4 && large_packet_stg3)) &&
                   (lower_padded_stg2 || framing_dsc_stg2)) begin
        pr_phyr_tlast_d    = 1'b1;
        tlast_on_mid_crc_d = 1'b0;
        packet_discontinue = (standard_dsc_case || framing_dsc_stg2 ||
                              stalled_discontinue || prx_cs_crc_check_fail[3]);
      // clean up after the last beat
      end else if (PR_phyr_tlast && PR_phyr_tvalid && !(set_eop_stg3 || eop_delay_stg3)) begin
        pr_phyr_tlast_d    = 1'b0;
        tlast_on_mid_crc_d = 1'b0;
        packet_discontinue = 1'b0;
      // discontinue due to destination (buffer), packet (stomp, lreq, etc), or error
      end else if (PR_phyr_tvalid && (standard_dsc_case || stalled_discontinue)) begin
        pr_phyr_tlast_d    = 1'b1;
        tlast_on_mid_crc_d = 1'b0;
        packet_discontinue = 1'b1;
      // lost link initialization, gracefully exit any packet transfer we're in the middle of
      end else if (!out_of_packet && !rt_stream_enable_stg2) begin
        pr_phyr_tlast_d    = 1'b1;
        tlast_on_mid_crc_d = 1'b0;
        packet_discontinue = 1'b1;
      // standard case -
      end else begin
        pr_phyr_tlast_d    = set_eop_stg3 || tvalid_delay;
        tlast_on_mid_crc_d = 1'b0;
        packet_discontinue = (set_eop_stg3 || tvalid_delay) &&
   //                          (standard_dsc_case || stalled_discontinue || (PR_phyr_tlast && PR_phyr_tuser[0])); // org logic
                             (standard_dsc_case || prx_in_recoverable_detect_delay || stalled_discontinue || (PR_phyr_tlast && PR_phyr_tuser[0]));
      end
    end else begin
      tlast_on_mid_crc_d = 1'b0;
      pr_phyr_tlast_d    = PR_phyr_tlast;
      packet_discontinue = PR_phyr_tuser[0];
    end
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      stalled_discontinue <= #TCQ 1'b0;
    //end else if ((PR_phyr_tvalid && BR_phyr_tready) || out_of_packet) begin
    end else if (out_of_packet) begin
      stalled_discontinue <= #TCQ 1'b0;
    end else begin
      stalled_discontinue <= #TCQ standard_dsc_case || (stalled_discontinue && !PR_phyr_tuser[0]);
    end
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PR_phyr_tlast     <= #TCQ 1'b0;
      tlast_on_mid_crc  <= #TCQ 1'b0;
      PR_phyr_tuser[0]  <= #TCQ 1'b0;
      large_packet_stg4 <= #TCQ 1'b0;
    end else begin
      PR_phyr_tlast     <= #TCQ pr_phyr_tlast_d;
      tlast_on_mid_crc  <= #TCQ tlast_on_mid_crc_d;
  //  PR_phyr_tuser[0]  <= #TCQ packet_discontinue; // org logic
      PR_phyr_tuser[0]  <= #TCQ pr_phyr_tlast_d ?
                                (packet_discontinue
                                             || PR_phyr_tuser[0]
                                             || prx_in_recoverable_detect_delay // CR# 849823
                                                 ) : 1'b0; // updated condition
      large_packet_stg4 <= #TCQ large_packet_stg3;
    end
  end


  // TSTRB generation -
  // the final byte enable is based on how much pad got added.
  // 32 bits of pad can be added to complete a packet.
  // 16 bits of pad can be added after the CRC.
  wire [3:0]   final_crc_loc       = (tvalid_delay && !out_of_packet) ? crc_loc_stg4 :
                                      single_cycle_stg3  ? crc_loc_stg2 : crc_loc_stg3;
  wire [3:0]   final_crc_loc_early = (tvalid_delay && !out_of_packet) ? crc_loc_stg3 : crc_loc_stg2;
  always @(posedge phy_clk) begin
    crc_loc_stg4 <= #TCQ crc_loc_stg3;
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PR_phyr_tkeep <= #TCQ 8'hFF;
    end else if (advance_condition
                 &&
                 pr_phyr_tlast_d
                ) begin
      // next three conditions are where the last beat contains no actual data.
      if (final_crc_loc_early == 4'h8 && !large_packet_stg3) begin
        PR_phyr_tkeep <= #TCQ 8'h7F;
      end else if (final_crc_loc_early == 4'h8 && large_packet_stg3 && lower_padded_stg2) begin
        PR_phyr_tkeep <= #TCQ 8'h1F;
      end else if (final_crc_loc_early == 4'h4 && large_packet_stg3 && lower_padded_stg2) begin
        PR_phyr_tkeep <= #TCQ 8'h7F;
      // last beat is where the mid crc would be
      end else if (mid_crc_loc_stg2 && framing_end_stg2) begin
        PR_phyr_tkeep <= #TCQ 8'h7F;
      end else begin
        case ({final_crc_loc, large_packet_stg3})
        5'b0001_0  : PR_phyr_tkeep <= #TCQ 8'h1F;
        5'b0001_1  : PR_phyr_tkeep <= #TCQ 8'h07;
        5'b0010_0  : PR_phyr_tkeep <= #TCQ 8'h07;
        5'b0010_1  : PR_phyr_tkeep <= #TCQ 8'h01;
        5'b0100_0  : PR_phyr_tkeep <= #TCQ 8'h01;
        5'b0100_1  : PR_phyr_tkeep <= #TCQ 8'h1F;
        default    : PR_phyr_tkeep <= #TCQ 8'hFF;
        endcase
      end
    end else begin
      PR_phyr_tkeep <= #TCQ 8'hFF;
    end
  end


  // TDATA generation -
  // byte shift and swizzle the data before going across AXI.
  assign PR_phyr_tdata = {phyr_tdata[7:0], phyr_tdata[15:8],  phyr_tdata[23:16], phyr_tdata[31:24],
                          phyr_tdata[39:32], phyr_tdata[47:40], phyr_tdata[55:48], phyr_tdata[63:56]};
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      phyr_tdata <= #TCQ 64'h0;
    end else if (advance_condition && !tvalid_delay) begin
      if (large_packet_stg3) begin // past the mid-crc
        phyr_tdata[63:24] <= #TCQ ordered_rx_data_stg3[39:0];
        phyr_tdata[23:0]  <= #TCQ ordered_rx_data_stg2[63:40];
      end else if (mid_crc_loc_stg2) begin // remove the mid-crc
        phyr_tdata[63:8]  <= #TCQ ordered_rx_data_stg3[55:0];
        phyr_tdata[7:0]   <= #TCQ ordered_rx_data_stg2[47:40];
      end else begin // anything before the mid-crc, only remove ackid
        phyr_tdata[63:8]  <= #TCQ ordered_rx_data_stg3[55:0];
        phyr_tdata[7:0]   <= #TCQ ordered_rx_data_stg2[63:56];
      end
    end
  end


  // TUSER generation - {1'b0, skip_crc, 3'h0, VC, CRF, src_dsc}
  // first 7 bits only need to be valid on the fist beat of a packet
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PR_phyr_tuser[7:1]  <= #TCQ 8'h0;
    end else if (advance_condition && !tvalid_delay) begin
      PR_phyr_tuser[7:1]  <= #TCQ {1'h0, SWITCH_MODE, 3'h0, vc_stg3, crf_stg3};
    end
  end


  // TVALID generation -
  always @(posedge phy_clk) begin
    if (phy_rst_q)
      out_of_packet <= #TCQ 1'b1;
    else if (PR_phyr_tvalid && BR_phyr_tready)
      out_of_packet <= #TCQ PR_phyr_tlast;
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PR_phyr_tvalid <= #TCQ 1'b0;
      tvalid_delay   <= #TCQ 1'b0;
    end else if (advance_condition) begin
      // special case #1:
      // swallow a packet that is being discontinued on or before the first beat
 //     if ((input_error_ns == IN_ERROR_RECOVERY) && !PR_phyr_tvalid && !(pr_phyr_tlast_d && !PR_phyr_tvalid))begin       // fix for CR 824332
 //     if ((input_error_cs == IN_ERROR_RECOVERY) && !PR_phyr_tvalid  && !PR_phyr_tlast && !pr_phyr_tlast_d)begin       // fix for CR 824332 // new addition
 //       PR_phyr_tvalid <= #TCQ 1'b0;
 //       tvalid_delay   <= #TCQ 1'b0;
//          end else if ((out_of_packet && !(PR_phyr_tvalid && BR_phyr_tready)) &&
          //end else if (((out_of_packet && !(PR_phyr_tvalid && BR_phyr_tready)) ||
      //     (PR_phyr_tvalid && BR_phyr_tready && PR_phyr_tlast)) &&
          if ((out_of_packet && !(PR_phyr_tvalid && BR_phyr_tready)) &&
           (standard_dsc_case || (!vc_stg3 && (!rt_stream_enable_stg3 || !rt_stream_enable_stg2)) ||
            ((crc_loc_stg2 == 4'h8) && (framing_dsc_stg2 || prx_cs_crc_check_fail[3])))) begin
        PR_phyr_tvalid <= #TCQ 1'b0;
        tvalid_delay   <= #TCQ 1'b0;
        end else if ((PR_phyr_tvalid && BR_phyr_tready) &&   // newly added logic RX fix                                    // fix for CR 822472
           ((prx_in_recoverable_detect_delay && !pr_phyr_tlast_d) || (!vc_stg3 && (!rt_stream_enable_stg3 || (!rt_stream_enable_stg2 && !pr_phyr_tlast_d))) ||
  //          ((crc_loc_stg2 == 4'h8) && (framing_dsc_stg2 || prx_cs_crc_check_fail[3])))) begin
            ((crc_loc_stg2 == 4'h8) && ((framing_dsc_stg3 && !pr_phyr_tlast_d) || prx_cs_crc_check_fail[3])))) begin   // 09_29(1)
        PR_phyr_tvalid <= #TCQ 1'b0; // newly added RC fix
        tvalid_delay   <= #TCQ 1'b0; // newly added RC fix
      // special case #2:
      // remove a final beat of a packet when it only contains crc.
      end else if (((crc_loc_stg3 == 4'h8) || (crc_loc_stg3 == 4'h4 && large_packet_stg4)) &&
                   !tvalid_delay && lower_padded_stg3 && !packet_discontinue) begin
        PR_phyr_tvalid <= #TCQ 1'b0;
        tvalid_delay   <= #TCQ 1'b0;
      // special case #3:
      // hold off tvalid when eop location causes a dead space
      end else if (eop_delay_stg3 && !pr_phyr_tlast_d) begin // added  && !pr_phyr_tlast_d, CR#825620
        PR_phyr_tvalid <= #TCQ 1'b0;
        tvalid_delay   <= #TCQ rt_stream_enable_stg3 && rt_stream_enable_stg2;
      // special case #4:
      // when the last beat is on the mid crc, kill a final, unneeded tvalid
      end else if (tlast_on_mid_crc) begin
        PR_phyr_tvalid <= #TCQ 1'b0;
        tvalid_delay   <= #TCQ 1'b0;
      // standard case
      end else begin
        //PR_phyr_tvalid <= #TCQ data_vld_stg3 || tvalid_delay || stalled_discontinue || pr_phyr_tlast_d;
        //PR_phyr_tvalid <= #TCQ data_vld_stg3 || tvalid_delay || pr_phyr_tlast_d;
        PR_phyr_tvalid <= #TCQ (
                                (data_vld_stg3 || tvalid_delay || pr_phyr_tlast_d)
                                &&
                                !(
                                                   (prx_in_recoverable_detect_delay && !pr_phyr_tlast_d)//CR# 851964
                                   &&
                                   !PR_phyr_tvalid
                                   &&
                                   !tvalid_delay
                                                 )
                                );    // fix for CR 821476, updated for RC fix
        tvalid_delay   <= #TCQ 1'b0;
      end
    end
  end


    // *- COVERAGE (cp_PR_eop_next_value)
    // See that EOP gets tagged with stage1 data

    // *- COVERAGE (cp_PR_eop_current_value)
    // See that EOP gets tagged with stage2 data

    // *- ASSERTION (ap_PR_src_dsc_on_first_beat)
    // src_dsc will never assert on the first cycle of a packet

  // }}} End of RX Buf Interface ----------

// }}} End Stage4 Pipeline ---------------

endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
//
// OLLM_RX_CS_DECODE
// Description:
// This module instantiates all the submodules of the OLLM RX design
//
// Hierarchy:
// PHY_TOP
//    |___OLLM_RX_TOP
//             |___OLLM_RX_CS_DECODE <-- this module
//             |_____OLLM_RX_DATAPATH
//             |_____OLLM_RX_ERR_DETECT
// ---------------------------------------------------------------------

`timescale 1ps/1ps

module srio_gen2_v4_1_16_ollm_rx_cs_decode
  #(
    parameter TCQ           = 100)  // in pS
   (
  // {{{ port declarations ----------------
    // clocks and resets and general signals
    input             phy_clk,                    // PHY interface clock
    input             phy_rst_q,                  // Reset for PHY clock Domain

    // OPLM Interface
    input      [63:0] PP_rx_data,                 // Receive data
    input      [7:0]  PP_rx_charisk,              // Indicates which bytes are K characters
    input      [1:0]  PP_rx_valid,                // Indicates valid words
    input             PP_idle2_selected,          // Indicates when an IDLE2 sequence is present
    input             PP_port_initialized,        // Indicates port is initialized
    input             PR_link_initialized,        // Indicates link is initialized

    // OPLM Interface
    output reg [63:0] PRD_rx_data,                // Receive data
    output reg [7:0]  PRD_rx_charisk,             // Indicates which bytes are K characters
    output reg [1:0]  PRD_rx_valid,               // Indicates valid words
    output reg        PRD_idle2_selected,         // Indicates when an IDLE2 sequence is present
    output reg [81:0] PRD_cs_decode,              // A whole series of control symbol decodes. See assignment
    output reg        idle2_sync_char_stg0
  // }}} ----------------------------------
   );

  // {{{ local parameters -----------------

  // Special Character decodes
  localparam [7:0] PD                    = 8'b011_11100; // K28.3
  localparam [7:0] SC                    = 8'b000_11100; // K28.0
  localparam [7:0] K_CHAR                = 8'b101_11100; // K28.5
  localparam [7:0] R_CHAR                = 8'b111_11101; // K29.7
  localparam [7:0] A_CHAR                = 8'b111_11011; // K27.7
  localparam [7:0] M_CHAR                = 8'b001_11100; // K28.1

  // Stype1 decodes
  localparam [2:0] C_SOP                 = 3'b000;
  localparam [2:0] C_STMP                = 3'b001;
  localparam [2:0] C_EOP                 = 3'b010;
  localparam [2:0] C_RFR                 = 3'b011;
  localparam [2:0] C_LREQ                = 3'b100;
  localparam [2:0] C_MCE                 = 3'b101;
  localparam [2:0] C_RSVD1               = 3'b110;
  localparam [2:0] C_NOP                 = 3'b111;

  // Stype0 decodes
  localparam [2:0] C_PA                  = 3'b000;
  localparam [2:0] C_PR                  = 3'b001;
  localparam [2:0] C_PNA                 = 3'b010;
  localparam [2:0] C_RSVD0               = 3'b011;
  localparam [2:0] C_STAT                = 3'b100;
  localparam [2:0] C_VSTAT               = 3'b101;
  localparam [2:0] C_LRESP               = 3'b110;
  localparam [2:0] C_IMP_DEF             = 3'b111;

  // CMD decodes
  localparam [2:0] C_LREQ_RST_DEV        = 3'b011; // sub-command for link request
  localparam [2:0] C_LREQ_IN_STAT        = 3'b100; // sub-command for link request

  // }}} End local parameters -------------


  // {{{ wire declarations ----------------
  // Prefix notation:
  // phy = phy clock domain
  // pr/PR = Physical Layer Receive
  // pt/PT = Physical Layer Transmit
  // pc/PC = Physical Layer Config
  // pp/PP = Physical Layer OPLM
  // br/BR = Buffer Layer Receive
  // prx   = Physical Layer Error Detection signals (Not 'pre' to avoid confusion)
  // _st*  = Pipeline Stage Number

  // - Data Parser
  reg   [1:0]            pd_flag;                  // Packet Delimiter Delimiter indication
  reg   [1:0]            sc_flag;                  // Control Symbol Delimiter indication
  wire  [2:0]            stype1_lower_bitsel;      // location of stype1 function in lower half
  wire  [2:0]            stype1_upper_bitsel;      // location of stype1 function in upper half
  wire  [2:0]            cmd_lower_bitsel;         // location of stype1 function in lower half
  wire  [2:0]            cmd_upper_bitsel;         // location of stype1 function in upper half
  wire  [2:0]            stype0_lower_bitsel;      // location of stype1 function in lower half
  wire  [2:0]            stype0_upper_bitsel;      // location of stype1 function in upper half
  wire  [5:0]            param0_lower_bitsel;      // location of parameter0 in the lower half
  wire  [5:0]            param0_upper_bitsel;      // location of parameter0 in the upper half
  wire  [5:0]            param1_lower_bitsel;      // location of parameter1 in the lower half
  wire  [5:0]            param1_upper_bitsel;      // location of parameter1 in the upper half

  // - Stype1 Decode
  reg   [1:0]            in_packet;                // indicates when the the data stream is part of a packet
  reg                    framing_start;            // used with in_packet to indicate the start of a packet
  reg                    framing_end;              // used with in_packet to indicate the end of a packet
  reg                    framing_dsc;              // used with in_packet to indicate a discontinued packet
  reg                    framing_dsc_delay;        // used with in_packet to indicate a discontinued packet
  wire  [1:0]            sop;                      // successful decode of SOP in either upper or lower
  wire  [1:0]            stomp;                    // successful decode of STOMP in either upper or lower
  wire  [1:0]            eop;                      // successful decode of EOP in either upper or lower
  wire  [1:0]            rfr;                      // successful decode of RFR in either upper or lower
  wire  [1:0]            lreq;                     // successful decode of LREQ in either upper or lower
  wire  [1:0]            lreq_rst_dev;             // successful decode of LREQ-rst-dev in either upper or lower
  wire  [1:0]            lreq_in_stat;             // successful decode of LREQ-in-stat in either upper or lower
  wire  [1:0]            mce;                      // successful decode of MCE in either upper or lower
  wire  [1:0]            s1rsvd;                   // successful decode of RSVD in either upper or lower
  wire  [1:0]            nop;                      // successful decode of NOP in either upper or lower

  // - Stype0 Decode
  wire  [5:0]            pa_ackid;                 // sampled from parameter0 - pa ackid
  wire  [5:0]            pr_ackid;                 // sampled from parameter0 - pr ackid
  wire  [5:0]            ackid_status;             // sampled from parameter0
  wire  [2:0]            vcid;                     // sampled from parameter0
  wire  [4:0]            port_status;              // sampled from parameter1
  wire  [5:0]            buf_status;               // sampled from parameter1
  wire  [4:0]            cause;                    // sampled from parameter1
  wire  [1:0]            pa;                       // successful decode of PA in either upper or lower
  wire  [1:0]            pr;                       // successful decode of PR in either upper or lower
  wire  [1:0]            pna;                      // successful decode of PNA in either upper or lower
  wire  [1:0]            s0rsvd;                   // successful decode of RSVD in either upper or lower
  wire  [1:0]            stat;                     // successful decode of STATUS in either upper or lower
  wire  [1:0]            vcstat;                   // successful decode of VC STATUS in either upper or lower
  wire  [1:0]            lresp;                    // successful decode of LRESP in either upper or lower
  wire  [1:0]            id;                       // successful decode of ID in either upper or lower

  // outgoing signal
  wire [81:0]            prd_cs_decode_d;          // unregistered bus of outgoing decodes. See assignment for mapping

  // common use signals
  reg pp_port_initialized_q;


  // }}} End wire declarations ------------


  // {{{ + Data Parser ----------------------
  // main interface to the OPLM. Register some stuff and create some
  // useful signals.

  always @(posedge phy_clk) begin
    pp_port_initialized_q   <= #TCQ PP_port_initialized;
  end

  // Generate the Packet Delimiter and Control Symbol signals.
  // They are seperate for error detection logic.
  wire [7:0] upper_delim_bitsel = PP_rx_data[63:56]; // only valid location for upper cs delimiter
  wire [7:0] lower_delim_bitsel = PP_rx_data[31:24]; // only valid location for lower cs delimiter
  wire [7:0] upper_extended_delim_bitsel = PP_rx_data[39:32]; // only valid location for upper cs delimiter
  wire [7:0] lower_extended_delim_bitsel = PP_rx_data[7:0]; // only valid location for lower cs delimiter
  always @* begin
    pd_flag = 2'h0;
    sc_flag = 2'h0;
    if (PP_rx_charisk[3] && pp_port_initialized_q) begin
      pd_flag[0] = lower_delim_bitsel == PD;
      sc_flag[0] = lower_delim_bitsel == SC;
    end
    if (PP_rx_charisk[7] && pp_port_initialized_q) begin
      pd_flag[1] = upper_delim_bitsel == PD;
      sc_flag[1] = upper_delim_bitsel == SC;
    end
  end

  // gather the bits used to decode stype1 functions.
  wire [2:0] short_stype1_lower_bitsel = PP_rx_data[10:8];  // location of stype1 for short/lower cs
  wire [2:0] long_stype1_lower_bitsel  = PP_rx_data[8:6];   // location of stype1 for long/lower cs
  wire [2:0] short_stype1_upper_bitsel = PP_rx_data[42:40]; // location of stype1 for short/upper cs
  wire [2:0] long_stype1_upper_bitsel  = PP_rx_data[40:38]; // location of stype1 for long/upper cs

  assign stype1_lower_bitsel = PRD_idle2_selected == 1 ? long_stype1_lower_bitsel: short_stype1_lower_bitsel;
  assign stype1_upper_bitsel = PRD_idle2_selected == 1 ? long_stype1_upper_bitsel: short_stype1_upper_bitsel;

  // gather the bits used to decode stype1 cmd.
  wire [2:0] short_cmd_lower_bitsel = PP_rx_data[7:5];   // location of cmd for short/lower cs
  wire [2:0] long_cmd_lower_bitsel  = PP_rx_data[5:3];   // location of cmd for long/lower cs
  wire [2:0] short_cmd_upper_bitsel = PP_rx_data[39:37]; // location of cmd for short/upper cs
  wire [2:0] long_cmd_upper_bitsel  = PP_rx_data[37:35]; // location of cmd for long/upper cs

  assign cmd_lower_bitsel = PRD_idle2_selected == 1 ? long_cmd_lower_bitsel: short_cmd_lower_bitsel;
  assign cmd_upper_bitsel = PRD_idle2_selected == 1 ? long_cmd_upper_bitsel: short_cmd_upper_bitsel;

  // gather the bits used to decode stype0 functions.
  wire [2:0] short_stype0_lower_bitsel = PP_rx_data[23:21]; // location of stype0 for short/lower cs
  wire [2:0] long_stype0_lower_bitsel  = PP_rx_data[23:21]; // location of stype0 for long/lower cs
  wire [2:0] short_stype0_upper_bitsel = PP_rx_data[55:53]; // location of stype0 for short/upper cs
  wire [2:0] long_stype0_upper_bitsel  = PP_rx_data[55:53]; // location of stype0 for long/upper cs

  assign stype0_lower_bitsel = PRD_idle2_selected == 1 ? long_stype0_lower_bitsel: short_stype0_lower_bitsel;
  assign stype0_upper_bitsel = PRD_idle2_selected == 1 ? long_stype0_upper_bitsel: short_stype0_upper_bitsel;

  // gather the bits used to decode parameter0.
  wire [5:0] short_param0_lower_bitsel = {1'b0, PP_rx_data[20:16]}; // location of parameter0 for short/lower cs
  wire [5:0] long_param0_lower_bitsel  = PP_rx_data[20:15];         // location of parameter0 for long/lower cs
  wire [5:0] short_param0_upper_bitsel = {1'b0, PP_rx_data[52:48]}; // location of parameter0 for short/upper cs
  wire [5:0] long_param0_upper_bitsel  = PP_rx_data[52:47];         // location of parameter0 for long/upper cs

  assign param0_lower_bitsel = PRD_idle2_selected == 1 ? long_param0_lower_bitsel: short_param0_lower_bitsel;
  assign param0_upper_bitsel = PRD_idle2_selected == 1 ? long_param0_upper_bitsel: short_param0_upper_bitsel;

  // gather the bits used to decode parameter1.
  wire [5:0] short_param1_lower_bitsel = {1'b0, PP_rx_data[15:11]}; // location of parameter1 for short/lower cs
  wire [5:0] long_param1_lower_bitsel  = PP_rx_data[14:9];          // location of parameter1 for long/lower cs
  wire [5:0] short_param1_upper_bitsel = {1'b0, PP_rx_data[47:43]}; // location of parameter1 for short/upper cs
  wire [5:0] long_param1_upper_bitsel  = PP_rx_data[46:41];         // location of parameter1 for long/upper cs

  assign param1_lower_bitsel = PRD_idle2_selected == 1 ? long_param1_lower_bitsel: short_param1_lower_bitsel;
  assign param1_upper_bitsel = PRD_idle2_selected == 1 ? long_param1_upper_bitsel: short_param1_upper_bitsel;


  // }}} End of Data Parser ---------------


  // {{{ + Stype1 Decode --------------------
  // all things related to the decode of Stype1 -
  // packet framing, stomps, link requests, multi-cast events
  reg [1:0] sop_q;
  reg       eop_q;
  reg       in_packet_q; // reduced from 1:0 to supress warnings
  reg [2:0] reset_device_cnt;

  // control symbol decode
  assign sop    = {(pd_flag[1] || sc_flag[1]) && stype1_upper_bitsel == C_SOP,
                   (pd_flag[0] || sc_flag[0]) && stype1_lower_bitsel == C_SOP};
  assign stomp  = {(pd_flag[1] || sc_flag[1]) && stype1_upper_bitsel == C_STMP,
                   (pd_flag[0] || sc_flag[0]) && stype1_lower_bitsel == C_STMP};
  assign eop    = {(pd_flag[1] || sc_flag[1]) && stype1_upper_bitsel == C_EOP,
                   (pd_flag[0] || sc_flag[0]) && stype1_lower_bitsel == C_EOP};
  assign rfr    = {(pd_flag[1] || sc_flag[1]) && stype1_upper_bitsel == C_RFR,
                   (pd_flag[0] || sc_flag[0]) && stype1_lower_bitsel == C_RFR};
  assign lreq   = {(pd_flag[1] || sc_flag[1]) && stype1_upper_bitsel == C_LREQ,
                   (pd_flag[0] || sc_flag[0]) && stype1_lower_bitsel == C_LREQ};
  assign mce    = {(pd_flag[1] || sc_flag[1]) && stype1_upper_bitsel == C_MCE,
                   (pd_flag[0] || sc_flag[0]) && stype1_lower_bitsel == C_MCE};
  assign s1rsvd = {sc_flag[1] && stype1_upper_bitsel == C_RSVD1,
                   sc_flag[0] && stype1_lower_bitsel == C_RSVD1};
  assign nop    = {sc_flag[1] && stype1_upper_bitsel == C_NOP,
                   sc_flag[0] && stype1_lower_bitsel == C_NOP};

  assign lreq_rst_dev = {lreq[1] && cmd_upper_bitsel == C_LREQ_RST_DEV,
                         lreq[0] && cmd_lower_bitsel == C_LREQ_RST_DEV};
  assign lreq_in_stat = {lreq[1] && cmd_upper_bitsel == C_LREQ_IN_STAT,
                         lreq[0] && cmd_lower_bitsel == C_LREQ_IN_STAT};


  // When determining the beginning of a packet, look for SOP one word
  // prior. When determining the close of a packet, look for any of the
  // ending delimiters on the same cycle. If neither of these occur,
  // take the previous value of the packet status.
  always @* begin
    if (sop_q[0] && !stomp[1])
      in_packet[1] = PR_link_initialized;
    else if (eop_q)
      in_packet[1] = 1'b0;
    else if ((lreq[1] || stomp[1]) && sop[0])// CR 825747
      in_packet[1] = 1'b0;                   // when BFM cancells packet (with stomp or lreq), dont send PNA   
    else
      in_packet[1] = in_packet_q;

    if (sop[1] && !stomp[0])
      in_packet[0] = PR_link_initialized;
    else if (eop[1] || stomp[1] || rfr[1] || lreq[1]) // any eop
      in_packet[0] = 1'b0;
    else
      in_packet[0] = in_packet[1];
  end

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      sop_q       <= #TCQ 0;
      eop_q       <= #TCQ 0;
      in_packet_q <= #TCQ 0;
    end else begin
      sop_q       <= #TCQ sop;
      eop_q       <= #TCQ eop[0] || stomp[0] || rfr[0] || lreq[0]; // any eop
      in_packet_q <= #TCQ in_packet[0];
    end
  end


  // Creation of the framing signals. These are single-cycle pulses
  // at the beginning, end, and whenever there is a discontinue.
  always @* begin
    if ((sop[1] && !stomp[0]) || (sop_q[0] && !stomp[1]))
      framing_start = 1'b1;
    else
      framing_start = 1'b0;

    if ((sop[1] || eop[1] || rfr[1] || (~|sop_q && lreq[1]) || (~|sop_q && stomp[1])) && in_packet[1])
      framing_end = 1'b1;
    else if ((sop[0] || eop[0] || rfr[0] || (!(sop[1] || sop_q[0]) && lreq[0]) ||
             (!(sop[1] || sop_q[0]) && stomp[0])) && in_packet[0])
      framing_end = 1'b1;
    else
      framing_end = framing_dsc_delay;

    if ((rfr[1] || (~|sop_q && lreq[1]) || (~|sop_q && stomp[1])) && in_packet[1])
      framing_dsc = 1'b1;
    else if ((rfr[0] || (!(sop[1] || sop_q[0]) && lreq[0]) ||
             (!(sop[1] || sop_q[0]) && stomp[0])) && in_packet[0])
      framing_dsc = 1'b1;
    else
      framing_dsc = framing_dsc_delay;
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      framing_dsc_delay <= #TCQ 1'b0;
    end else if ((sop_q[1] && (stomp[1] || lreq[1])) || (sop_q[0] && (stomp[0] || lreq[0]))) begin
      framing_dsc_delay <= #TCQ 1'b1;
    end else begin
      framing_dsc_delay <= #TCQ 1'b0;
    end
  end

//----- below code checks the IDLE2 sync sequence CR #820674 -------------------
  wire [7:0] idle2_m_char;
  assign idle2_m_char[7] = (|sop_q || |in_packet) ? ((PP_rx_data[63:56] == M_CHAR) && PP_rx_charisk[7]) : 1'b0;
  assign idle2_m_char[6] = (|sop_q || |in_packet) ? ((PP_rx_data[55:48] == M_CHAR) && PP_rx_charisk[6]) : 1'b0;
  assign idle2_m_char[5] = (|sop_q || |in_packet) ? ((PP_rx_data[47:40] == M_CHAR) && PP_rx_charisk[5]) : 1'b0;
  assign idle2_m_char[4] = (|sop_q || |in_packet) ? ((PP_rx_data[39:32] == M_CHAR) && PP_rx_charisk[4]) : 1'b0;

  assign idle2_m_char[3] = (|sop_q || |in_packet) ? ((PP_rx_data[31:24] == M_CHAR) && PP_rx_charisk[3]) : 1'b0;
  assign idle2_m_char[2] = (|sop_q || |in_packet) ? ((PP_rx_data[23:16] == M_CHAR) && PP_rx_charisk[2]) : 1'b0;
  assign idle2_m_char[1] = (|sop_q || |in_packet) ? ((PP_rx_data[15:8]  == M_CHAR) && PP_rx_charisk[1]) : 1'b0;
  assign idle2_m_char[0] = (|sop_q || |in_packet) ? ((PP_rx_data[7:0]   == M_CHAR) && PP_rx_charisk[0]) : 1'b0;

  reg idle2_sync_char;
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
        idle2_sync_char_stg0 <= 1'b0;
    end else begin
        idle2_sync_char_stg0 <= idle2_sync_char;
    end
  end

  always @* begin : check_idle2_sync_char
      if (!PP_port_initialized) begin
        idle2_sync_char     = 1'b0;
      end else if (!PP_idle2_selected) begin
        idle2_sync_char     = 1'b0;
      end else begin
        if (|idle2_m_char     // if M char is present on any of the lanes
            &&
            !(|lreq)
            &&
            |in_packet        // packet has been started
            ) begin
          idle2_sync_char = 1'b1;
        end else begin
          idle2_sync_char = idle2_sync_char_stg0   // The asserted signal will de-assert
                            &&                // when LREQ is received
                            !(|lreq);
        end
      end
  end
//----- code which checks the IDLE2 sync sequence CR #820674 ends --------------

  // }}} End of Stype1 Decode -------------


  // {{{ + Stype0 Decode --------------------

  reg   [5:0]            pa_ackid_q;
  reg   [5:0]            pr_ackid_q;
  reg   [5:0]            ackid_status_q;
  reg   [2:0]            vcid_q;
  reg   [5:0]            buf_status_q;
  reg   [4:0]            cause_q;
  reg   [4:0]            port_status_q;

  // control symbol decode
  assign pa     = {(pd_flag[1] || sc_flag[1]) && stype0_upper_bitsel == C_PA,
                   (pd_flag[0] || sc_flag[0]) && stype0_lower_bitsel == C_PA};
  assign pr     = {(pd_flag[1] || sc_flag[1]) && stype0_upper_bitsel == C_PR,
                   (pd_flag[0] || sc_flag[0]) && stype0_lower_bitsel == C_PR};
  assign pna    = {(pd_flag[1] || sc_flag[1]) && stype0_upper_bitsel == C_PNA,
                   (pd_flag[0] || sc_flag[0]) && stype0_lower_bitsel == C_PNA};
  assign s0rsvd = {(pd_flag[1] || sc_flag[1]) && stype0_upper_bitsel == C_RSVD0,
                   (pd_flag[0] || sc_flag[0]) && stype0_lower_bitsel == C_RSVD0};
  assign stat   = {(pd_flag[1] || sc_flag[1]) && stype0_upper_bitsel == C_STAT,
                   (pd_flag[0] || sc_flag[0]) && stype0_lower_bitsel == C_STAT};
  assign vcstat = {(pd_flag[1] || sc_flag[1]) && stype0_upper_bitsel == C_VSTAT,
                   (pd_flag[0] || sc_flag[0]) && stype0_lower_bitsel == C_VSTAT};
  assign lresp  = {(pd_flag[1] || sc_flag[1]) && stype0_upper_bitsel == C_LRESP,
                   (pd_flag[0] || sc_flag[0]) && stype0_lower_bitsel == C_LRESP};
  assign id     = {(pd_flag[1] || sc_flag[1]) && stype0_upper_bitsel == C_IMP_DEF,
                   (pd_flag[0] || sc_flag[0]) && stype0_lower_bitsel == C_IMP_DEF};


  // Parameter0 updates - packet_ackid
  assign pa_ackid      = pa[0] ? param0_lower_bitsel :
                         pa[1] ? param0_upper_bitsel :
                         pa_ackid_q;
  assign pr_ackid      = pr[0] ? param0_lower_bitsel :
                         pr[1] ? param0_upper_bitsel :
                         pr_ackid_q;

  // Parameter0 updates - ackid_status
  // NOTE: ackid_status is also passed with a status control symbol.
  // It is not as reliable as the value we're keeping internally
  // and not collected here.
  assign ackid_status      = lresp[0] ? param0_lower_bitsel :
                             lresp[1] ? param0_upper_bitsel :
                             ackid_status_q;

  // Parameter0 updates - vcid
  assign vcid      = vcstat[0] ? param0_lower_bitsel[2:0] :
                     vcstat[1] ? param0_upper_bitsel[2:0] :
                     vcid_q;


  // Parameter1 updates - buf_status
  // NOTE: buf_status is also passed with a VC_status control symbol.
  // This is not the same buffer status as the others, and
  // not collected here.
  assign buf_status      =  (pa[0] || pr[0] || stat[0]) ? param1_lower_bitsel :
                            (pa[1] || pr[1] || stat[1]) ? param1_upper_bitsel :
                            buf_status_q;

  // Parameter1 updates - cause
  // NOTE: Cause field isn't used for anything at the moment.
  assign cause      = pna[0] ? param1_lower_bitsel[4:0] :
                      pna[1] ? param1_upper_bitsel[4:0] :
                      cause_q;

  // Parameter1 updates - port_status
  assign port_status      = lresp[0] ? param1_lower_bitsel[4:0] :
                            lresp[1] ? param1_upper_bitsel[4:0] :
                            port_status_q;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      pa_ackid_q     <= #TCQ 0;
      pr_ackid_q     <= #TCQ 0;
      ackid_status_q <= #TCQ 0;
      vcid_q         <= #TCQ 0;
      buf_status_q   <= #TCQ 0;
      cause_q        <= #TCQ 0;
      port_status_q  <= #TCQ 0;
    end else begin
      pa_ackid_q     <= #TCQ pa_ackid;
      pr_ackid_q     <= #TCQ pr_ackid;
      ackid_status_q <= #TCQ ackid_status;
      vcid_q         <= #TCQ vcid;
      buf_status_q   <= #TCQ buf_status;
      cause_q        <= #TCQ cause;
      port_status_q  <= #TCQ port_status;
    end
  end

  // }}} End of Stype0 Decode -------------


  // {{{ + Final Register -------------------
  assign prd_cs_decode_d = {
                            // Data parser [81:78]
                            pd_flag,       // [81:80]
                            sc_flag,       // [79:78]

                            // Stype1 [77:53]
                            in_packet,     // [77:76]
                            framing_start, // [75]
                            framing_end,   // [74]
                            framing_dsc,   // [73]
                            sop,           // [72:71]
                            stomp,         // [70:69]
                            eop,           // [68:67]
                            rfr,           // [66:65]
                            lreq,          // [64:63]
                            lreq_rst_dev,  // [62:61]
                            lreq_in_stat,  // [60:59]
                            mce,           // [58:57]
                            s1rsvd,        // [56:55]
                            nop,           // [54:53]

                            // Stype0 [52:0]
                            pa_ackid,      // [52:47]
                            pr_ackid,      // [46:41]
                            ackid_status,  // [40:35]
                            vcid,          // [34:32]
                            port_status,   // [31:27]
                            buf_status,    // [26:21]
                            cause,         // [20:16]
                            pa,            // [15:14]
                            pr,            // [13:12]
                            pna,           // [11:10]
                            s0rsvd,        // [9:8]
                            stat,          // [7:6]
                            vcstat,        // [5:4]
                            lresp,         // [3:2]
                            id};           // [1:0]


  always @(posedge phy_clk) begin
    PRD_rx_data        <= #TCQ PP_rx_data;
    PRD_idle2_selected <= #TCQ PP_idle2_selected;
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PRD_rx_charisk     <= #TCQ 0;
      PRD_rx_valid       <= #TCQ 0;
      PRD_cs_decode      <= #TCQ 0;
    end else begin
      PRD_rx_charisk     <= #TCQ PP_rx_charisk;
      PRD_rx_valid       <= #TCQ PP_rx_valid;
      PRD_cs_decode      <= #TCQ prd_cs_decode_d;
    end
  end

  // }}} End of Final Register ------------


endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/phy/ollm_rx/srio_gen2_v4_1_16_ollm_rx_err_detect.v#2 $
//----------------------------------------------------------------------
//
// OLLM_RX_ERR_DETECT
// Description:
// This module instantiates all of the error detection logic for the
// OLLM_RX
//
// Hierarchy:
// PHY_TOP
//    |___OLLM_RX_TOP
//             |_____OLLM_RX_DATAPATH
//             |_____OLLM_RX_ERR_DETECT <-- this module
// ---------------------------------------------------------------------

`timescale 1ps/1ps

module srio_gen2_v4_1_16_ollm_rx_err_detect
  #(
    parameter TCQ           = 100,  // in pS
    parameter IDLE1         = 1,    // Include the IDLE1 sequence {0, 1}
    parameter IDLE2         = 0,    // Include the IDLE2 sequence {0, 1}
    parameter MODE_XG       = 5,    // Line rates {1/1.25, 2/2.5, 3/3.125, 5/5, 6/6.25}
    parameter VC            = 0,    // Highest number VC supported {0, 1}
    parameter SWITCH_MODE   = 0,    // If the core is generated with Switch Mode Support {0, 1}
    parameter RETRY         = 1,    // Includes Retry protocol {0, 1}
    parameter LINK_REQUESTS = 3,    // Additional link requests to send prior to port_error {0, 1, 2, 3, 4, 5, 6, 7}
    parameter LINK_WIDTH    = 1)          // Number of GT lanes to use {1, 2, 4}

   (
  // {{{ port declarations ----------------
    // clocks and resets and general signals
    input             phy_clk,                    // PHY interface clock
    input             phy_rst_q,                  // Reset for PHY clock Domain
    input             log_clk,                    // LOG interface clock
    input             log_rst_q,                  // Reset for LOG clock Domain
    input             gt_pcs_clk,                 // GT interface clock

    // external inputs
    input      [63:0] PRD_rx_data,                // Receive data
    input      [7:0]  PRD_rx_charisk,             // Indicates which bytes are K characters
    input             PRD_idle2_selected,         // Indicates when an IDLE2 sequence is present
    input      [LINK_WIDTH*4-1:0] PP_gt_decode_error,       // INVALID on GT RX (notintable or disperr)
    input             PP_mode_1x,                 // Indicates core has trained down to 1x // updated to fix CR# 835498

    input             PR_phyr_tvalid,             // Valid data indicator
    input             BR_phyr_tready,             // Destination Ready
    input             PR_phyr_tlast,              // Last DW of incoming packet
    input      [7:0]  PR_phyr_tuser,              // {1'h0, skip_crc, 3'h0, VC, CRF, src_dsc} AXI Compliance Pad
    input      [4:0]  PR_port_stat,               // Current port status
    input             PR_port_stat_ok,            // Port Status is OK
    input             PR_link_initialized,        // Indicates we are ready to transmit data
    input             PT_sample_next_fm,          // Indicates to the ollm rx to sample the next fm

    input      [5:0]  BR_phy_buf_stat,            // Buffer status from the RX Buffer
    input      [5:0]  PC_next_rcvd_pkt,           // Load value for Next Expected packet
    input      [5:0]  PC_last_ack,                // Load value for phy_last_ack when Pload_ackids is asserted
    input             PC_load_ackids,             // Loads next_rcvd_pkt with CFG provided alternatives
    input             PC_load_nextpkt,            // Load next_rcvd_pkt with CFG value
    input             PC_send_lreq,               // Send a Link Request Input Status CS
    input       [2:0] PC_lreq_cmd,                // Command information for PC_send_lreq
    input      [23:0] PC_link_timeout,            // Time-out value for packet acknowledgement
    input             PC_input_maint_only,        // Only maintenance traffic is allowed
    input      [5:0]  PT_phy_next_fm,             // Next Packet's Ack ID
    input             PR_output_error_stop,       // OLLM RX is currently in Output Error Stopped State
    input             PR_output_retry_stop,       // OLLM RX is currently in Output Retry Stopped State
    input             PR_input_status_good,       // OLLM RX is currently in Input Waiting for Event State
    input             PR_send_pna,                // Send a PNA control symbol
    input             PR_send_lreq,               // Send a LREQ control symbol
    input             PT_lreq_sent,               // Sent Link Request
    input      [5:0]  PR_ackid_status,            // sampled from parameter0
    input             err_recovery,
    input             carryover_stg2,
    input      [1:0]  data_vld_stg0_d,            // Delayed data valid to identify charisk


    // external outputs
    output reg [4:0]  PRX_cause,                  // Last cause for a PNA to send
    output     [5:0]  PRX_phy_last_ack,           // Last PA received by the PHY core
    output     [5:0]  PRX_last_good_pkt,          // Last PA to send
    output     [5:0]  PRX_next_rcvd_pkt,          // Next expected packet AckID
    output reg        PRX_phy_rcvd_mce,           // MCE control symbol received
    output    [31:0]  prx_debug,                  // debug signals for error detection module



    // internal datapath inputs
    // stage 0
    input      [1:0]  pd_flag_stg0,               // Packet Delimiter Delimiter indication
    input      [1:0]  sc_flag_stg0,               // Control Symbol Delimiter indication
    input      [1:0]  in_packet_stg0,             // Indicates when in or out of a packet
    input      [1:0]  sop,                        // successful decode of SOP in either upper or lower
    input      [1:0]  stomp,                      // successful decode of STOMP in either upper or lower
    input      [1:0]  eop,                        // successful decode of EOP in either upper or lower
    input      [1:0]  rfr,                        // successful decode of RFR in either upper or lower
    input      [1:0]  lreq,                       // successful decode of LREQ in either upper or lower
    input      [1:0]  stat,                       // successful decode of STAT in either upper or lower
    input      [1:0]  mce,                        // successful decode of MCE in either upper or lower

    // stage 1
    input      [63:0] masked_rx_data_stg1,        // Receive data, masked AckID for CRC check
    input      [63:0] ordered_rx_data_stg1,       // Receive data
    input             data_vld_stg1,              // data valid window
    input             data_stream_enable_stg1,    // stream enable for both RT and CT
    input             pp_out_of_sync_stg1,        // Scrambler is out of sync
    input             pp_port_initialized_stg1,   // Indicates port is initialized
    input      [3:0]  crc_loc_stg1,               // one-hot location for the CRC
    input             mid_crc_loc_stg1,           // Beat identifier for the mid CRC
    input             beat_count_q_is_10,         // Just might be the location of the mid-crc
    input             framing_end_stg1,           // indicates the end of a packet
    input             framing_start_stg1,         // indicates the start of a packet
    input             framing_dsc_stg1,           // used with in_packet to indicate a discontinued packet
    input             upper_valid_stg1,           // Data valid signal after reordering for AXI
    input             lower_valid_stg1,           // Data valid signal after reordering for AXI
    input             lower_padded_stg1,          // when 1, the lower word is pad at the end of a packet
    input             first_beat_stg1,            // first beat of a packet
    input             stomp_detect_stg1,          // Stomp control symbol received
    input             lresp_detect_stg2,          // Link-Response identifier
    input      [1:0]  pa_detect_stg1,             // Packet-Ack identifier
    input      [1:0]  pa_detect_stg0,             // 2/5/2015
    input             pr_detect_stg1,             // Packet-Retry identifier
    input             rfr_detect_stg1,            // Restart-from-Retry identifier
    input             lreq_detect_stg1,           // Link-Request identifier
    input      [1:0]  lreq_in_stat_detect_stg1,   // Link-Request detection - in stat
    input      [5:0]  pa_ackid_stg1,              // sampled from parameter0 - pa ackid
    input      [5:0]  pr_ackid_stg1,              // sampled from parameter0 - pr ackid
    input      [1:0]  expected_ackid_coef_stg1,   // when two PAs, value of 2, otherwise 1

    // stage 2
    input             framing_end_stg2,           // indicates the end of a packet
    input             framing_start_stg2,         // used with in_packet to indicate the start of a packet
    input       [3:0] crc_loc_stg2,               // one-hot location for the CRC
    input             mid_crc_loc_stg2,           // Beat identifier for the mid CRC
    input             rt_stream_enable_stg2,      // Used to enable the stream for RT
    input             dest_dsc_stg2,              // Determination for destination discontinue

    // outputs consumed by datapath
    output            prx_out_fatal_detect,       // Output fatal error condition discovered
    output reg        prx_force_send_lreq,        // Forces the OLLM TX to send a LREQ
    output            prx_out_recoverable_detect, // Output recoverable error condition discovered
    output            prx_in_recoverable_detect,  // Input recoverable error condition discovered
    output            prx_in_retry_detect,        // Retry condition discovered
    output reg  [3:0] prx_cs_crc_check_fail,      // used to generate cs_crc_in_error_cond
    output reg        prx_cs_in_error_cond,       // control symbol error condition detected
    output reg        prx_rcvd_bad_status,        // Asserts when there is an error in status
    input             idle2_sync_char_stg0,       // added to fix idle2 based CR #820674
    input             in_retry_stopped_state,     // added to indicate the input retry stopped state
    output            control_sym_in_error_cond_cmb, //
    input             not_in_retry_stopped_state, // used to check the next state in CR 825487 fixes
    output            idle_seq_in_error_cond_cmb, // added to pass the combo error to datapath satemachine
    output            lreq_pd_error,
    input  [1:0]      lreq_reset_dev,             // detects the LREQ+RST
    input             in_error_stopped_state,     // added to ignore any errors when in error stopped state,
                                                  // CR# 837481

    output            idle2_7_4_beat_err_cmb      // CR# 849824
  // }}} ----------------------------------
   );

  // {{{ local parameters -----------------

  // Special Character decodes
  localparam [7:0] PD                    = 8'b011_11100; // K28.3
  localparam [7:0] SC                    = 8'b000_11100; // K28.0
  localparam [7:0] K_CHAR                = 8'b101_11100; // K28.5
  localparam [7:0] R_CHAR                = 8'b111_11101; // K29.7
  localparam [7:0] A_CHAR                = 8'b111_11011; // K27.7
  localparam [7:0] M_CHAR                = 8'b001_11100; // K28.1

  // For encoding the Cause field
  localparam [4:0] C_UNEXPECTED_ACKID    = 5'b00001;
  localparam [4:0] C_BAD_CS_CRC          = 5'b00010;
  localparam [4:0] C_NON_MAINTENANCE     = 5'b00011;
  localparam [4:0] C_BAD_PACKET_CRC      = 5'b00100;
  localparam [4:0] C_INVALID_CHAR        = 5'b00101;
  localparam [4:0] C_RESOURCE_RETRY      = 5'b00110;
  localparam [4:0] C_LOSS_OF_SYNC        = 5'b00111;

  // FTYPE decode
  localparam [3:0] FTYPE_MAINT           = 4'b1000;

  // Based on MODE_XG, determine the upper bit of the SRL
  localparam       N_CNT_MAX = MODE_XG == 6 ? 31 :
                               MODE_XG == 5 ? 31 :
                               MODE_XG == 3 ? 15 :
                               MODE_XG == 2 ? 15 :
                               MODE_XG == 1 ?  7 :
                                               7;

  // Port Status
  localparam [4:0] PORT_STAT_ERROR       = 5'b00010;
  localparam [4:0] PORT_STAT_RETRY_STOP  = 5'b00100;
  localparam [4:0] PORT_STAT_ERROR_STOP  = 5'b00101;
  localparam [4:0] PORT_STAT_OK          = 5'b10000;

  // }}} End local parameters -------------


  // {{{ wire declarations ----------------

  // commonly used signals
  reg  [5:0]        prx_phy_last_ack_int;         // last_ack value before masking the upper bit
  reg               prx_in_recoverable_detect_q;  // Input recoverable error condition discovered
  wire              ok_ackid;                     // when 1, received ackid falls within a valid range in error
  wire [5:0]        expected_ackid;               // phy_last_ack + 1
  wire [5:0]        masked_expected_ackid;        // masked upper bit of above when in IDLE1
  reg               prx_in_retry_detect_q;        // registered retry detection
  wire              first_valid_beat_stg1;        // asserted on the very first beat of a packet
  reg  [1:0]        pd_flag_stg1;                 // packet delimiter
  reg  [1:0]        pd_flag_stg2;                 // packet delimiter
  reg  [1:0]        sc_flag_stg1;                 // packet delimiter - registered
  reg               cfg_requested_lresp;          // asserts when the user requested a lresp through registers
  reg  [3:0]        prx_cs_crc_check_fail_q;      // used to generate cs_crc_in_error_cond
  reg  [1:0]        pa_detect_stg2;
  reg  [1:0]        pa_detect_stg3;
  reg  [1:0]        bad_delimiter_stg1;           // packet is using a wrong delimiter
  reg  [1:0]        bad_delimiter_stg2;           // packet is using a wrong delimiter
  reg               pr_output_error_stop_q;
  reg               pr_output_retry_stop_q;

  // output fatal errors
  reg               link_timer_fatal_cond;        // any type of link timer output fatal error
  reg  [2:0]        overall_fatal_count;          // used for when the counter must expire multiple times
  reg               control_sym_fatal_cond;       // any type of control symbol output fatal error

  // output recoverable errors
  reg               link_timer_out_error_cond;    // any type of link timer output recoverable error
  wire              control_sym_out_error_cond;   // any type of control symbol output recoverable error
  reg [3:1]         control_sym_out_error_cond_d; // any type of control symbol output recoverable error

  // input recoverable errors
  reg               control_sym_in_error_cond;    // any type of control symbol input recoverable error
  reg [6:1]         control_sym_in_error_cond_d;  // bitwise selection of error condition
  reg               control_sym_in_error_straddle;// control symbol error straddles beat boundary
  reg               control_sym_in_error_straddle_d; // straddled across beat boundaries
  reg               idle_seq_in_error_cond;       // any type of IDLE sequence input recoverable error
  reg               packet_in_error_cond;         // any type of packet input recoverable error
  wire              crc_in_error_cond;            // any type of CRC input recoverable error
  wire                 pk_crc_in_error_cond;      // packet-only CRC error, subset of crc_in_error_cond
  reg                  cs_crc_in_error_cond;      // cs-only CRC error, subset of crc_in_error_cond
  reg                  cs_crc_in_error_cond_mod;  // modification of above to assert for a sorter pulse
  reg                  cs_crc_in_error_cond_mod_q;// modification of above to assert for a sorter pulse
  reg               ignore_pk_crc;                // When set, ignore packet crc errors due to other complications
  reg               prx_cs_crc_check_fail_early;  // used to generate cs_crc_in_error_cond
  reg               ackid_in_error_cond;          // any type of AckID input recoverable error
  reg               ackid_in_error_cond_q;        // any type of AckID input recoverable error
  reg               other_in_error_cond;          // other types of error conditions
  reg                  loss_of_sync;              // loss of sync only, subset of other_in_error_cond
  reg                  rcvd_non_maint_packet;     // non-maint packet, subset of other_in_error_cond
  wire              invalid_char_in_sync_seq;     // added to detect the invalid character in the sync sequence
  reg               idle2_sync_char_stg1;
  reg               idle2_sync_char_stg2;         // added 2 stage delay to fix the CR# 847695
  // input retry conditions
  reg               control_sym_retry_cond;       // any type of control symbol input recoverable error
  reg               control_sym_retry_cond_d;     // early version of above
  reg               rx_buf_retry_cond;            // any type of Buffer input retry
  wire              rx_buf_retry_cond_d;          // early of above
  wire              control_sym_in_error_cond_dd_cmb; // 2/5/2015
  reg [6:1]         control_sym_in_error_cond_dd = 6'h0; // unregistered control symbol error detection
  
  reg [7:0] PRD_rx_charisk_reg;
  reg [7:0] PRD_rx_charisk_reg2;

  reg       sc_pd_mismatch_stg1;
  reg      idle2_7_4_beat_err;
  reg      idle2_3_0_beat_err;
  reg       idle2_7_4_beat_err_reg;
  reg       idle2_3_0_beat_err_reg;

  // error detection logic signals
  (* shreg_extract = "yes" *)
  reg [N_CNT_MAX:0] n_counter = 15;               // SRL-based counter, translates link rate to duration
  reg [23:0]        link_timer;                   // link timer, designed to timeout between 3 and 6 seconds
  wire              link_timer_enable;            // allows the larger timer to incrment
  reg               link_timer_enable_q;          // allows the larger timer to incrment
  reg               framing_dsc_stg1_delay;       // Delayed framing disconnect

  // }}} End wire declarations ------------
  reg [3:0]         rx_charisk_stg1;
  reg [1:0]         lreq_rst_dev_detect_stg1; // 
  reg               lreq_rst_dev_detect_stg2; // 
  wire              control_sym_in_error_cond_dd_ORed; // 
  // {{{ prx_debug assignment --------------

// newly added functionality to detect the invalid characters duing the sync sequence,
// During sync sequence,when there are no PD or SC detected by the core and when charisk shows asserted, its
// and invalid error.
assign invalid_char_in_sync_seq = !(|sc_flag_stg0 || |pd_flag_stg0) // during sync sequence, when there are no SC or 
                                  &&				    // PD detected, but charisk is detected for
				  idle2_sync_char_stg1              // invalid SC/PD places, then generate an error
				  &&                                // CR# 847695
                                  (PRD_rx_charisk[7] && PRD_rx_charisk[0]);



  assign prx_debug = {
                      19'h0,
                      framing_dsc_stg1,                  // 1
                      framing_end_stg1,                  // 1
                      framing_start_stg1,                // 1
                      |in_packet_stg0,                   // 1
                      prx_in_recoverable_detect,         // 1
                      prx_in_retry_detect,               // 1
                      prx_out_recoverable_detect,        // 1
                      prx_out_fatal_detect,              // 1
                      PRX_cause                          // 5
                      };

  // }}} -----------------------------------

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
        idle2_sync_char_stg1 <= 1'b0;
	    idle2_sync_char_stg2 <= 1'b0;
    end else begin
        idle2_sync_char_stg1 <= idle2_sync_char_stg0;
        idle2_sync_char_stg2 <= idle2_sync_char_stg1 && !(|lreq);// added extra 2 staged delay
    end
  end
  // {{{ Commonly Used Signals ------------
  assign first_valid_beat_stg1 = first_beat_stg1 && data_vld_stg1 && data_stream_enable_stg1;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      pd_flag_stg1                <= #TCQ 2'b0;
      pd_flag_stg2                <= #TCQ 2'b0;
      sc_flag_stg1                <= #TCQ 2'b0;
      prx_in_recoverable_detect_q <= #TCQ 1'b0;
      pr_output_error_stop_q      <= #TCQ 1'b0;
      pr_output_retry_stop_q      <= #TCQ 1'b0;
      lreq_rst_dev_detect_stg1    <= #TCQ 2'h0;// 
      lreq_rst_dev_detect_stg2    <= #TCQ 1'b0;// 
    end else begin
      pd_flag_stg1                <= #TCQ pd_flag_stg0;
      pd_flag_stg2                <= #TCQ pd_flag_stg1;
      sc_flag_stg1                <= #TCQ sc_flag_stg0;
      prx_in_recoverable_detect_q <= #TCQ prx_in_recoverable_detect;
      pr_output_error_stop_q      <= #TCQ PR_output_error_stop;
      pr_output_retry_stop_q      <= #TCQ PR_output_retry_stop;
      lreq_rst_dev_detect_stg1    <= #TCQ |lreq_reset_dev && idle2_sync_char_stg1;//
      lreq_rst_dev_detect_stg2    <= #TCQ lreq_rst_dev_detect_stg1 && PRD_idle2_selected;// 
    end
  end

  // register the MultiCast Event. OLLM doesn't use this, only forwards it on.
  reg [1:0] mce_q;
  reg       mce_qq;
  reg       phy_rcvd_mce;
  reg [1:0] phy_rcvd_mce_sync;
  reg       phy_rcvd_mce_sync_q;
  reg       phy_rcvd_mce_sync_qq;
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      phy_rcvd_mce <= #TCQ 1'b0;
      mce_q        <= #TCQ 2'b00;
      mce_qq       <= #TCQ 1'b0;
    end else if (PR_link_initialized) begin
      mce_q        <= #TCQ mce;

      mce_qq       <= #TCQ !prx_cs_crc_check_fail[2] && !control_sym_in_error_cond_d[3] && !control_sym_in_error_cond_d[1] &&   // fix for CR 838089
                           ((mce_q[0] && !prx_cs_crc_check_fail[1] && !bad_delimiter_stg2[0]) ||
                           (mce_q[1] && !prx_cs_crc_check_fail[0] && !bad_delimiter_stg2[1]));

      phy_rcvd_mce <= #TCQ mce_qq && !prx_cs_crc_check_fail[3] && !control_sym_in_error_straddle;
    end
  end
  always @(posedge log_clk or posedge phy_rcvd_mce) begin
    if (phy_rcvd_mce) begin
      phy_rcvd_mce_sync <= #TCQ 2'b11;
    end else begin
      phy_rcvd_mce_sync <= #TCQ {phy_rcvd_mce_sync[0], 1'b0};
    end
  end
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      phy_rcvd_mce_sync_q  <= #TCQ 1'b0;
      phy_rcvd_mce_sync_qq <= #TCQ 1'b0;
      PRX_phy_rcvd_mce     <= #TCQ 1'b0;
    end else begin
      phy_rcvd_mce_sync_q  <= #TCQ |phy_rcvd_mce_sync;
      phy_rcvd_mce_sync_qq <= #TCQ phy_rcvd_mce_sync_q;
      PRX_phy_rcvd_mce     <= #TCQ !phy_rcvd_mce_sync_qq && phy_rcvd_mce_sync_q;
    end
  end

  // }}} End Commonly Used Signals --------

  reg gt_decode_error_pcs_clk_stg1;
  reg gt_decode_error_pcs_clk_stg2;

  (* ASYNC_REG = "TRUE" *)
  reg gt_decode_error_phy_clk_stg1;
  (* ASYNC_REG = "TRUE" *)
  reg gt_decode_error_phy_clk_stg2;

  always @(posedge gt_pcs_clk) begin // updated to fix CR# 835498
        gt_decode_error_pcs_clk_stg1 <= #TCQ pp_port_initialized_stg1 ?
                                        (PP_mode_1x ? |PP_gt_decode_error[3:0] : |PP_gt_decode_error)
                                        :
                                        1'b0 ;
        gt_decode_error_pcs_clk_stg2 <= #TCQ gt_decode_error_pcs_clk_stg1;
     end

  // updated to fix CR# 835498
  wire gt_decode_error = (pp_port_initialized_stg1 ? (PP_mode_1x ? |PP_gt_decode_error[3:0] :|PP_gt_decode_error) : 1'b0)
                         || gt_decode_error_pcs_clk_stg1 || gt_decode_error_pcs_clk_stg2;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
        gt_decode_error_phy_clk_stg1 <= #TCQ 1'b0;
        gt_decode_error_phy_clk_stg2 <= #TCQ 1'b0;
      end else begin
        gt_decode_error_phy_clk_stg1 <= #TCQ gt_decode_error;
        gt_decode_error_phy_clk_stg2 <= #TCQ gt_decode_error_phy_clk_stg1;
      end
    end

  // {{{ Final error and signal creation --

  // Error types
  assign prx_out_fatal_detect       = link_timer_fatal_cond || control_sym_fatal_cond;
  assign prx_out_recoverable_detect = link_timer_out_error_cond || control_sym_out_error_cond;
  assign prx_in_recoverable_detect  = control_sym_in_error_cond 
                                      || idle_seq_in_error_cond 
				                      || packet_in_error_cond 
				                      || crc_in_error_cond 
				                      || prx_cs_crc_check_fail_q[3] 
				                      || ackid_in_error_cond_q 
				                      || other_in_error_cond 
				                      || gt_decode_error_phy_clk_stg2
				                      || invalid_char_in_sync_seq;// added to fix the CR# 847695
  assign prx_in_retry_detect        = control_sym_retry_cond
                                      ||
                                      rx_buf_retry_cond
                                      ||
                                      lreq_rst_dev_detect_stg2
                                      ; // 

  always @(posedge phy_clk) begin
    if (phy_rst_q)
      prx_in_retry_detect_q <= #TCQ 1'b0;
    else
      prx_in_retry_detect_q <= #TCQ prx_in_retry_detect;
  end


  // Generate the Cause field for outgoing PNAs
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PRX_cause <= #TCQ 5'b11111;
    end else if (!PR_send_pna
                 &&
                 (
                   (
                     prx_in_recoverable_detect
                     &&
                     !prx_in_recoverable_detect_q
                   )
                   ||
                   (
                     prx_in_retry_detect
                     &&
                     !RETRY
                   )
                 )
                 ) begin
      casex (
      {(control_sym_in_error_cond 
        || 
	    packet_in_error_cond 
	    || 
	    gt_decode_error_phy_clk_stg2 
	    || 
	    invalid_char_in_sync_seq // added to detect the invalid characters in sync sequence for IDLE2, CR# 847695
       ),
       ackid_in_error_cond_q,
       rcvd_non_maint_packet,
       (prx_cs_crc_check_fail_q[3] || cs_crc_in_error_cond), // //CR# 835364 is fixed, removed _mod_q condition
       (pk_crc_in_error_cond && !ignore_pk_crc && PR_port_stat_ok),
       rx_buf_retry_cond,
       loss_of_sync}
       )
      7'b1xxxxxx : PRX_cause <= #TCQ C_INVALID_CHAR;
      7'b01xxxxx : PRX_cause <= #TCQ C_UNEXPECTED_ACKID;
      7'b001xxxx : PRX_cause <= #TCQ C_NON_MAINTENANCE;
      7'b0001xxx : PRX_cause <= #TCQ C_BAD_CS_CRC;
      7'b00001xx : PRX_cause <= #TCQ C_BAD_PACKET_CRC;
      7'b000001x : PRX_cause <= #TCQ C_RESOURCE_RETRY;
      7'b0000001 : PRX_cause <= #TCQ C_LOSS_OF_SYNC;
      default    : PRX_cause <= #TCQ 5'b11111;
      endcase
    end
  end

//--------------------------------------------------------------------------------
  `ifdef SIMULATION

    reg [25*8-1:0] prx_cause_string = "NONE";

    always @* begin
      //PRX_cause
      case (PRX_cause)
        5'b00001            : prx_cause_string = "C_UNEXPECTED_ACKID ";
        5'b00010            : prx_cause_string = "C_BAD_CS_CRC       ";
        5'b00011            : prx_cause_string = "C_NON_MAINTENANCE  ";
        5'b00100            : prx_cause_string = "C_BAD_PACKET_CRC   ";
        5'b00101            : prx_cause_string = "C_INVALID_CHAR     ";
        5'b00110            : prx_cause_string = "C_RESOURCE_RETRY   ";
        5'b00111            : prx_cause_string = "C_LOSS_OF_SYNC     ";
        default             : prx_cause_string = "NONE               ";
      endcase
     end
  `endif
//--------------------------------------------------------------------------------

  // Generate the expected phy_last_ack, output phy_last_ack when expected matches received
  reg  [5:0] prx_phy_last_ack_full;
  reg  [5:0] prx_phy_last_ack_full_q;


  // Generate phy_last_ack
  // IPCV - PRX_phy_last_ack[5] has a 2:1 mux when in IDLE2 and isn't directly registered
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      prx_phy_last_ack_full <= #TCQ 6'h3F;
    end else if (PC_load_ackids) begin
      prx_phy_last_ack_full <= #TCQ {PRD_idle2_selected & PC_last_ack[5], PC_last_ack[4:0]};
    end else if (PR_link_initialized && lresp_detect_stg2 && !prx_cs_crc_check_fail[3] && ok_ackid) begin
      prx_phy_last_ack_full <= #TCQ PR_ackid_status - 1;
    end else if (PR_link_initialized && |pa_detect_stg2 && !PRD_idle2_selected) begin
      prx_phy_last_ack_full <= #TCQ prx_phy_last_ack_int;
    // special consideration must be made for packets that straddle across beat boundaries.
    end else if (PR_link_initialized && PRD_idle2_selected) begin
      if (pa_detect_stg2[0] && !control_sym_out_error_cond && prx_cs_crc_check_fail[3]) begin
        prx_phy_last_ack_full <= #TCQ  prx_phy_last_ack_full_q;
      end else if (|pa_detect_stg3) begin
        prx_phy_last_ack_full <= #TCQ prx_phy_last_ack_int;
      end
    end
  end
  assign PRX_phy_last_ack = PRD_idle2_selected ? prx_phy_last_ack_full : {1'b0, prx_phy_last_ack_full[4:0]};

  assign     expected_ackid        = prx_phy_last_ack_int + expected_ackid_coef_stg1;
  assign     masked_expected_ackid = {expected_ackid[5] && PRD_idle2_selected, expected_ackid[4:0]};
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      pa_detect_stg2          <= #TCQ 2'b0;
      pa_detect_stg3          <= #TCQ 2'b0;
      prx_phy_last_ack_full_q <= #TCQ 6'h3F;
    end else begin
      pa_detect_stg2          <= #TCQ pa_detect_stg1;
      pa_detect_stg3          <= #TCQ pa_detect_stg2;
      if (!(pa_detect_stg2[0] && PRD_idle2_selected &&
          !control_sym_out_error_cond && prx_cs_crc_check_fail[3])) begin
        prx_phy_last_ack_full_q <= #TCQ prx_phy_last_ack_int;
      end
    end
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      prx_phy_last_ack_int <= #TCQ 6'h3F;
    end else if (PC_load_ackids) begin
      prx_phy_last_ack_int <= #TCQ {PRD_idle2_selected & PC_last_ack[5], PC_last_ack[4:0]};
    // special case - if there was a crc error on an IDLE2 control symbol that straddles across beats,
    // revert the internal count value to the last known good value.
    // Why not only change it when you know it's good? Because by the time we know it's good,
    // another ack might arrive and we'll consider it to be wrong.
    end else if (pa_detect_stg2[0]
                 &&
                 PRD_idle2_selected
                 &&
                 !control_sym_out_error_cond
                 &&
                 prx_cs_crc_check_fail[3]
                 ) begin
      prx_phy_last_ack_int <= #TCQ prx_phy_last_ack_full_q;

    end else if (pa_detect_stg1[0]
                 &&
                 !prx_cs_crc_check_fail[1]
                 &&
                 !control_sym_in_error_cond_d[3]
                 &&
                 !((control_sym_in_error_cond_d[1] && !(idle2_7_4_beat_err_reg && PRD_idle2_selected))// CR #849076
                    ||
		    (control_sym_in_error_cond_dd[1] && idle2_7_4_beat_err && PRD_idle2_selected) // CR 849822
		 )
                 &&
                 !bad_delimiter_stg2[0]
                 &&
                 !(pa_detect_stg1[1] && prx_cs_crc_check_fail[0])
                 &&
                 !control_sym_out_error_cond_d[1]
                 &&
                 !PR_output_error_stop
                 ) begin
      prx_phy_last_ack_int <= #TCQ pa_ackid_stg1;
    end else if (pa_detect_stg1[1]
                 &&
                 !control_sym_in_error_cond_d[3]
                 &
                 !(control_sym_in_error_cond_d[1] && !(idle2_7_4_beat_err_reg && PRD_idle2_selected))//CR #849076
                 &&
                 !bad_delimiter_stg2[1]
                 &&
                 !prx_cs_crc_check_fail[0]
                 &&
                 !prx_cs_crc_check_fail[2]
                 &&
                 !control_sym_out_error_cond_d[1]
                 &&
                 !PR_output_error_stop
                 ) begin
      prx_phy_last_ack_int <= #TCQ prx_phy_last_ack_int + 1; // do not use pa_ackid_stg1 incase of b2b PAs, w/crc err
    end else if (lresp_detect_stg2
                 &&
                 !prx_cs_crc_check_fail[3]
                 &&
                 ok_ackid) begin
      prx_phy_last_ack_int <= #TCQ PR_ackid_status - 1;
    end
  end

    // *- COVERAGE (cp_PRX_cause_enumerate)
    // Observe all valid values for PR_cause

    // *- ASSERTION (ap_PRX_cause_illegal)
    // PR_cause will never be Reserved

    // *- COVERAGE (cp_PRX_b2b_pa_with_proper_ackid)
    // Observe back to back PAs with the proper ackids

    // *- ASSERTION (cp_PRX_last_ack_invalid_incr)
    // PRX_phy_last_ack never increments by more than 1 or 2 outside of a rewind


  // }}} End Final error creation ---------


  // {{{ classes of error detections ------

  // {{{ + Link Timer ---------------------
  // Checks being performed:
  // Out Fatal Error
  // 1) Link-Request/Link-Response handshake timeout
  // Out Recoverable Error
  // 1) No acknowledgement on a sent packet


  // Infer the SRL -
  // This free-running counter should take advantage of the SRL architecture
  // and is intended to make it so that the overall counter expires
  // somewhere between 3 and 6 seconds, regardless of the link rate.
  // gt_pcs_clk frequency | N counter length
  // 62.5 MHz         | 32
  // 125 MHz          | 64
  // 156.25 MHz       | 64
  // 250 MHz          | 128
  // 312.5 MHz        | 128
  assign link_timer_enable = n_counter[N_CNT_MAX];
  always @(posedge phy_clk) begin
    link_timer_enable_q <= #TCQ link_timer_enable;
  end
  always @(posedge gt_pcs_clk) begin
    n_counter <= #TCQ {n_counter[N_CNT_MAX-1:0], n_counter[N_CNT_MAX]};
  end

  // Create the 24-bit counter -
  // We could use either gt_pcs_clk or phy_clk, since they are related
  // by frequency AND the clock enable (from the SRL) beats at
  // a normalized pace, regardless of lane count and link rate.
  // This counter is used for both fatal and non-fatal error detection.
  // Clear on -
  // 1) transition between error/retry/normal modes (fatal detect)
  // 2) no outstanding packets (recoverable detect)
  // 3) packet acknowledgement (recoverable detect)
  wire [5:0] phy_last_ack_plus_1 = PRX_phy_last_ack + 6'h01;
  reg        hold_link_timer;
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      link_timer      <= #TCQ 24'h0;
      hold_link_timer <= #TCQ 1'b0;
    end else if (hold_link_timer) begin
      link_timer      <= #TCQ 24'h0;
      hold_link_timer <= #TCQ !PT_lreq_sent;
    end else if ((PR_output_error_stop && !pr_output_error_stop_q) ||
                 (PR_output_retry_stop && !pr_output_retry_stop_q) || PR_send_lreq ||
                 (lresp_detect_stg2 && !prx_cs_crc_check_fail[3])) begin // 
      link_timer      <= #TCQ 24'h0;
    end else if (!PR_output_error_stop &&  PRD_idle2_selected &&
                 (PT_phy_next_fm == phy_last_ack_plus_1)) begin // 
      link_timer      <= #TCQ 24'h0;
    end else if (!PR_output_error_stop && !PRD_idle2_selected &&
                 (PT_phy_next_fm[4:0] == phy_last_ack_plus_1[4:0])) begin // 
      link_timer      <= #TCQ 24'h0;
    end else if (!PR_output_error_stop && (|pa_detect_stg1)) begin // 
      link_timer      <= #TCQ 24'h0;
    end else if ((link_timer >= PC_link_timeout) && overall_fatal_count < LINK_REQUESTS) begin
      link_timer      <= #TCQ 24'h0;
      hold_link_timer <= #TCQ !PT_lreq_sent;
    end else if ((link_timer_enable && !link_timer_enable_q) && (PC_link_timeout > link_timer)) begin
      link_timer      <= #TCQ link_timer + 1;
    end
  end


  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      overall_fatal_count       <= #TCQ 3'h0;
      prx_force_send_lreq       <= #TCQ 1'b0;
    end else if (!PR_output_error_stop) begin
      overall_fatal_count       <= #TCQ 3'h0;
      prx_force_send_lreq       <= #TCQ 1'b0;
    end else if ((link_timer >= PC_link_timeout) && overall_fatal_count < LINK_REQUESTS) begin
      overall_fatal_count       <= #TCQ overall_fatal_count + 1;
      prx_force_send_lreq       <= #TCQ 1'b1;
    end else begin
      prx_force_send_lreq       <= #TCQ 1'b0;
    end
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      link_timer_fatal_cond     <= #TCQ 1'b0;
      link_timer_out_error_cond <= #TCQ 1'b0;
    end else begin
      link_timer_fatal_cond     <= #TCQ (link_timer >= PC_link_timeout) && PR_output_error_stop &&
                                        !link_timer_out_error_cond && overall_fatal_count >= LINK_REQUESTS;
      link_timer_out_error_cond <= #TCQ (link_timer >= PC_link_timeout) && !PR_output_error_stop;
    end
  end


    // *- ASSERTION (ap_PRX_link_timer_behavior)
    // Link timer should not expire if no data is sent after recovering from an Output Error or Retry

    // *- COVERAGE (cp_PRX_cross_pa_timeout)
    // Observe a link timeout on a packet acknowledgment event crossed with all speeds

    // *- COVERAGE (cp_PRX_cross_lreq_timeout)
    // Observe a timeout on a Link-Request/Link-Response handshake crossed with all speeds

  // }}} End of Link Timer ----------------


  // {{{ + Control Symbol Error Detection -
  // Checks being performed:
  // Out Fatal Error
  //   1) Link Response with unexpected AckID
  // Out Recoverable Error
  //   1) Packet-Acknowledge with unexpected AckID
  //   2) Packet Retry on an unexpected AckID
  //   3) Link Response when no Link Request was sent
  // In Recoverable Error
  //   1a) Long control symbol that does not have the correct (or not at all) end delimiter
  //   1b) Long control symbol that does not have a beginning delimiter
  //   2) Control symbol that uses the wrong delimiter
  //   3) Control symbol with invalid or non-data character
  //   4) Restart-from-Retry when not expecting one
  //   5) Packet-Retry when in multi-VC mode
  //   6) End-of-Packet when not in packet
  // In Retry Condition
  //   1) Receipt of a Stomp control symbol


  // The acceptable values of AckID fall between last_ack and next_fm, not including next_fm
  // Also check to see if next_fm has wrapped under but last_ack hasn't yet.
  reg [5:0]  pt_phy_next_fm_copy;
  reg        ackid_status_less_than_next_fm;
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      pt_phy_next_fm_copy            <= #TCQ 0;
    end else if (!prx_out_recoverable_detect && !pr_output_error_stop_q) begin
      pt_phy_next_fm_copy    <= #TCQ PT_phy_next_fm;
    end else if (PT_sample_next_fm) begin
      pt_phy_next_fm_copy    <= #TCQ PT_phy_next_fm;
    end
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      ackid_status_less_than_next_fm <= #TCQ 1'b1;
    end else begin
      ackid_status_less_than_next_fm <= #TCQ PR_ackid_status <= pt_phy_next_fm_copy;
    end
  end
  assign ok_ackid = (pt_phy_next_fm_copy > PRX_phy_last_ack) ?
                     (PR_ackid_status > PRX_phy_last_ack) && ackid_status_less_than_next_fm :
                     (PR_ackid_status > PRX_phy_last_ack) || ackid_status_less_than_next_fm;


  // Out Fatal Error Detect -
  // 1) Link Response with an unexpected AckID
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      control_sym_fatal_cond <= #TCQ 1'b0;
    end else if (!pp_port_initialized_stg1) begin
      control_sym_fatal_cond <= #TCQ 1'b0;
    end else if (lresp_detect_stg2 && !prx_cs_crc_check_fail[3]) begin
      control_sym_fatal_cond <= #TCQ !ok_ackid;
    end else begin
      control_sym_fatal_cond <= #TCQ 1'b0;
    end
  end


  // Out Recoverable Error -

  // 1) Packet-Ack with an unexpected AckID
  always @* begin
    // miscompare when there is no crc error or control symbol error
    if (|pa_detect_stg1 && (pa_ackid_stg1 != masked_expected_ackid) &&
        ~|prx_cs_crc_check_fail[2:0] && !prx_cs_in_error_cond) begin
      control_sym_out_error_cond_d[1] = 1'b1;
    // b2b straddled pa, where the first one had a crc error
    end else if (|pa_detect_stg1 && |pa_detect_stg2 && prx_cs_crc_check_fail[3]) begin
      control_sym_out_error_cond_d[1] = 1'b1;
    // b2b same cycle pa, where the first one had a crc error
    end else if (&pa_detect_stg1 && prx_cs_crc_check_fail[0]) begin
      control_sym_out_error_cond_d[1] = 1'b1;
    // PA when there are no free ids to ack
    end else if (|pa_detect_stg1 && !prx_cs_in_error_cond &&
                 ({PT_phy_next_fm[5] && PRD_idle2_selected, PT_phy_next_fm[4:0]} ==
                  {prx_phy_last_ack_int[5] && PRD_idle2_selected, prx_phy_last_ack_int[4:0]} + 6'h1)) begin
      control_sym_out_error_cond_d[1] = 1'b1;
    end else begin
      control_sym_out_error_cond_d[1] = 1'b0;
    end
  end

  // 2) Packet Retry on an unexpected AckID
  // Must be last_ack + 1
  reg pr_detect_stg1_q = 0;
  always @(posedge phy_clk) begin
    pr_detect_stg1_q <= #TCQ pr_detect_stg1 && ~|prx_cs_crc_check_fail[2:0];
  end
  always @* begin
    if (pr_detect_stg1_q && !prx_cs_crc_check_fail[3])
      control_sym_out_error_cond_d[2] = pr_ackid_stg1 != masked_expected_ackid;
    else
      control_sym_out_error_cond_d[2] = 1'b0;
  end

  // 3) Link Response when no Link Request was sent
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      cfg_requested_lresp <= #TCQ 1'b0;
    end else if (PC_send_lreq && PC_lreq_cmd == 3'b100) begin
      cfg_requested_lresp <= #TCQ 1'b1;
    end else if (lresp_detect_stg2 && !prx_cs_crc_check_fail[3]) begin
      cfg_requested_lresp <= #TCQ 1'b0;
    end
  end
  always @* begin
    if (lresp_detect_stg2 && !prx_cs_crc_check_fail[3])
      control_sym_out_error_cond_d[3] = !(PR_output_error_stop || cfg_requested_lresp);
    else
      control_sym_out_error_cond_d[3] = 1'b0;
  end

  reg control_sym_out_error_cond_raw;
  always @(posedge phy_clk) begin
    if (phy_rst_q)
      control_sym_out_error_cond_raw <= #TCQ 1'b0;
    else
      control_sym_out_error_cond_raw <= #TCQ (|control_sym_out_error_cond_d && !control_sym_in_error_straddle_d);
  end

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PRD_rx_charisk_reg  <= #TCQ 8'b0;
      PRD_rx_charisk_reg2 <= #TCQ 8'b0;
    end else begin
      PRD_rx_charisk_reg <= #TCQ PRD_rx_charisk;// 
      PRD_rx_charisk_reg2 <= #TCQ PRD_rx_charisk_reg;// 
    end 
  end
  

  wire idle2_control_sym_error_cond;
  assign idle2_control_sym_error_cond = (
                                        PRD_idle2_selected 
                                        && 
                                        control_sym_in_error_cond_dd_cmb 
                                        && 
                                        pa_detect_stg0[0] 
                                        &&
                                        PRD_rx_charisk[3]
                                        &&
                                        !(
                                          (PRD_rx_charisk[4] )//
                                          ||
                                          (PRD_rx_charisk_reg[3]  )//
                                         )
                                      )
                                      ||
                                      (
                                        PRD_idle2_selected 
                                        && 
                                        control_sym_in_error_cond_dd_cmb 
                                        && 
                                        pa_detect_stg0[1] 
                                        &&
                                        (PRD_rx_charisk[0] 
                                        || 
                                        PRD_rx_charisk[7])
                                      );

  assign control_sym_out_error_cond = (control_sym_out_error_cond_raw && !prx_cs_crc_check_fail[3])
                                      ;


  // In Recoverable Error -
  // NOTE - extra register added on this category of error to improve timing
  //reg [6:1] control_sym_in_error_cond_dd = 6'h0; // unregistered control symbol error detection

  // 1a) Long control symbol that does not have the correct (or not at all) end delimiter
  // 1b) Long control symbol that does not have a beginning delimiter
  reg       lower_delimiter_q;
  reg [7:0] lower_delimiter_data_q;
  reg       control_sym_compare;
  always @(posedge phy_clk) begin
    lower_delimiter_q      <= #TCQ (pd_flag_stg0[0] || sc_flag_stg0[0]);
    lower_delimiter_data_q <= #TCQ PRD_rx_data[31:24];
    control_sym_compare    <= #TCQ !(PRD_rx_data[63:56] == PRD_rx_data[7:0]) || !PRD_rx_charisk[0];
  end

reg [3:0] control_sym_in_error_cond_dd_4_bit;

  always @* begin
    // 1a)
    // long control symbol is completely represented in a single 64-bits

    control_sym_in_error_straddle_d = 1'b0;
    idle2_7_4_beat_err = 1'b0;
    idle2_3_0_beat_err = 1'b0;

    control_sym_in_error_cond_dd_4_bit = 4'b0;
    if (
        PRD_idle2_selected 
        && 
	    (pd_flag_stg0[1] || sc_flag_stg0[1]) 
	    &&
        (!(PRD_rx_data[63:56] == PRD_rx_data[7:0]) || !PRD_rx_charisk[0] || !PRD_rx_charisk[7])
	    ) begin

      control_sym_in_error_cond_dd_4_bit[0] = 1'b1;
    end
    // 1a)
    // long control symbol is straddled over two beats
    if (PRD_idle2_selected 
        && 
	    lower_delimiter_q 
	    &&
        (!(lower_delimiter_data_q == PRD_rx_data[39:32]) || !PRD_rx_charisk[4])
	) begin

      control_sym_in_error_cond_dd_4_bit[1] = 1'b1;
      control_sym_in_error_straddle_d = 1'b1;
      idle2_7_4_beat_err = 1'b1;
    end
    // 1b)
    // long control symbol is completely represented in a single 64-bits
    if (PRD_idle2_selected 
        && 
	    PRD_rx_charisk[3:0] == 4'b0001 
	    &&
        ((PRD_rx_data[7:0] == PD) || (PRD_rx_data[7:0] == SC)) 
	    && 
	    (!pd_flag_stg0[1] && !sc_flag_stg0[1])
	    ) begin

      control_sym_in_error_cond_dd_4_bit[2] = 1'b1;
    end
    // 1b)
    // long control symbol is straddled over two beats
    if (PRD_idle2_selected 
        && 
	    PRD_rx_charisk[7:4] == 4'b0001 
	    &&
        ((PRD_rx_data[39:32] == PD) || (PRD_rx_data[39:32] == SC)) 
	    && 
	    !lower_delimiter_q
	    ) begin

      control_sym_in_error_cond_dd_4_bit[3] = 1'b1;
      control_sym_in_error_straddle_d = 1'b1;
      idle2_7_4_beat_err = 1'b1;
    end
  end

always @* begin
   control_sym_in_error_cond_dd[1] = |control_sym_in_error_cond_dd_4_bit;
end

always @(posedge phy_clk) begin
  if (phy_rst_q) begin
      idle2_7_4_beat_err_reg <= #TCQ 1'b0;
  end else begin
      idle2_7_4_beat_err_reg <= #TCQ idle2_7_4_beat_err;
  end
end

assign idle2_7_4_beat_err_cmb = idle2_7_4_beat_err; // CR# 849824, 2/23/2015

//__ start of new logic addition _______________________________________________
// 11/27/2014, CR #834779
//__ below logic is added to check the PD errors for LREQ. In such cases core should
//__  stop sending the lresp from the input error statemachine in the datapath file.
//__ the below logic targets to check the LREQ PD errors in IDLE2 cases, in all beat conditions
//__ mentioned above for control_sym_in_error_cond_dd[1] cases

reg lreq_combined_stg0;

always @(posedge phy_clk) begin:reg_and_combine_lreq
  if (phy_rst_q) begin
      lreq_combined_stg0 <= #TCQ 1'b0;
  end else if (lreq_combined_stg0) begin
      lreq_combined_stg0 <= #TCQ 1'b0;
  end else begin
      lreq_combined_stg0 <= #TCQ |(lreq);
  end
end

wire lreq_pd_error_cmb;
assign lreq_pd_error_cmb = PRD_idle2_selected?
                           (control_sym_in_error_cond_d[1] && lreq_combined_stg0)
                           :
                           control_sym_in_error_cond_dd[1] && (|lreq || lreq_combined_stg0); // 


reg lreq_pd_error_stg0;
always @(posedge phy_clk) begin:register_lreq_pd_error
  if (phy_rst_q) begin
      lreq_pd_error_stg0 <= #TCQ 1'b0;
  end else if (lreq_pd_error_cmb) begin
      lreq_pd_error_stg0 <= #TCQ 1'b1;
  end else if (|lreq && !control_sym_in_error_cond_dd[1]) begin
      lreq_pd_error_stg0 <= #TCQ 1'b0;
  end
end
//___ ___|-|_______ lreq_pd_error_cmb
//___ _____|------- lreq_pd_error_stg0
assign lreq_pd_error = lreq_pd_error_stg0 || lreq_pd_error_cmb;
//___ ___|-|_______ lreq_pd_error_cmb
//___ _____|------- lreq_pd_error_stg0
//___ ___|--------- lreq_pd_error -- goes to Input error recovery state machine

//__ end of new logic addition _________________________________________________


  // 2) Control symbol that uses the wrong delimiter

//______________Start : To fix the CR# 825487 below logic is added _____________
//__When the IDLE1 core is in Retry stopped state, the only way to come out is
//__to provide the RFR.Below logic update checks the PD errors in RFR generation

reg sop_asserted;
reg sop_asserted_stg0;

always @* begin :idle1_sop_in_retry_stopped_state
    if (!PRD_idle2_selected && in_retry_stopped_state) begin
          if (sop[1] && !(|rfr) && !sop_asserted_stg0) begin
              sop_asserted = 1'b1;
          end else if (sop[0] && !(|rfr) && !sop_asserted_stg0) begin
              sop_asserted = 1'b1;
          end else if (|eop || |rfr) begin
              sop_asserted = 1'b0;
          end else begin
              sop_asserted = sop_asserted_stg0;
          end
    end else begin
        sop_asserted = 1'b0;
    end
end

always @(posedge phy_clk) begin
  sop_asserted_stg0 <= #TCQ sop_asserted;
end

reg rfr_pd_1_error;
reg rfr_pd_0_error;

// use below code for future updates if any 
// always @* begin :idle1_chk_pd_errors_for_rfr
//    if (
//        (sop_asserted_stg0 && (sop[0])
//        &&
//         (
//          ((PRD_rx_data[63:56] == PD) && (PRD_rx_data[42:40] == 3'b011) && !PRD_rx_charisk[7])
//          ||
//          (!(PRD_rx_data[63:56] == PD) && (PRD_rx_data[42:40] == 3'b011) && PRD_rx_charisk[7])
//         )
//         )
//        ) begin
//        rfr_pd_1_error = !not_in_retry_stopped_state; // 1'b1;
//    end else if (
//        (sop_asserted_stg0 && (eop[1] || sop[1])
//         &&
//         (
//          (((PRD_rx_data[31:24] == SC)) && (PRD_rx_data[10:8] == 3'b011) && !PRD_rx_charisk[3])
//          ||
//          (!((PRD_rx_data[31:24] == SC)) && (PRD_rx_data[10:8] == 3'b011) && PRD_rx_charisk[3])
//         )
//        )
//        )
//       begin
//        rfr_pd_0_error = !not_in_retry_stopped_state; // 1'b1;
//    end else begin
//        rfr_pd_1_error = 1'b0;
//        rfr_pd_0_error = 1'b0;
//    end
// end
 always @* begin :idle1_chk_pd_errors_for_rfr1
    if (
        (
         sop_asserted_stg0
         &&
         (sop[0])
         &&
         (
          ((PRD_rx_data[63:56] == PD) && (PRD_rx_data[42:40] == 3'b011) && !PRD_rx_charisk[7])
          ||
          (!(PRD_rx_data[63:56] == PD) && (PRD_rx_data[42:40] == 3'b011) && PRD_rx_charisk[7])
         )
        )
       ) begin
        rfr_pd_1_error = !not_in_retry_stopped_state; // 
    end else begin
        rfr_pd_1_error = 1'b0;
    end
 end

 always @* begin :idle1_chk_pd_errors_for_rfr0
    if (
        (
         sop_asserted_stg0
         &&
         (eop[1] || sop[1])
         &&
         (
          (((PRD_rx_data[31:24] == SC)) && (PRD_rx_data[10:8] == 3'b011) && !PRD_rx_charisk[3])
          ||
          (!((PRD_rx_data[31:24] == SC)) && (PRD_rx_data[10:8] == 3'b011) && PRD_rx_charisk[3])
         )
        )
       )
       begin
        rfr_pd_0_error = !not_in_retry_stopped_state; // 
    end else begin
        rfr_pd_0_error = 1'b0;
    end
 end

//______________End : To fix the CR# 825487 above logic is added in bad_delimiter_stg1 bits __

  always @* begin
    bad_delimiter_stg1[1] = (
                             (pd_flag_stg0[1] ^ (sop[1] || stomp[1] || eop[1]))
                             &&
                             !(rfr[1] || lreq[1])
                            )
                             ||
                             (pd_flag_stg0[1] && mce[1])
                             ||                       // Added to fix the CR 824965
                             (                        //
                              pd_flag_stg0[1]         // RFR should not be at
                              &&                      // packet delimter when
                              in_retry_stopped_state  // NOt in the packet and
                              &&                      // core is retry stopped state
                              rfr[1]                  //
                              &&                      //
                              !in_packet_stg0[1]      //
                              )                       //
                            //  ||                      // Added to fix the CR
                            //  rfr_pd_1_error          // 825487, idle1 case
                             ;

    bad_delimiter_stg1[0] = (
                             (pd_flag_stg0[0] ^ (sop[0] || stomp[0] || eop[0]))
                             &&
                             !(rfr[0] || lreq[0])
                            )
                             ||
                             (pd_flag_stg0[0] && mce[0])
                             ||                          //
                             (                           //
                              pd_flag_stg0[0]            // Added to fix the CR 824965
                              &&                         // RFR should not be at
                              in_retry_stopped_state     // packet delimter when
                              &&                         // NOt in the packet and
                              rfr[0]                     // core is retry stopped state
                              &&                         //
                              !in_packet_stg0[0]         //
                              )
                        //      ||                         // Added to fix the CR
                        //      rfr_pd_0_error             // 825487, idle1 case
                             ;
  end

  always @(posedge phy_clk) begin
    bad_delimiter_stg2 <= bad_delimiter_stg1;
  end
  always @* begin
    control_sym_in_error_cond_dd[2] = |bad_delimiter_stg1;
  end

  // 3) Control symbol with invalid or non-data character
  always @* begin
    // short in upper and/or lower
    if (!PRD_idle2_selected && (|pd_flag_stg0 || |sc_flag_stg0))
      control_sym_in_error_cond_dd[3] = ((pd_flag_stg0[1] || sc_flag_stg0[1]) && |PRD_rx_charisk[6:4]) ||
                                             ((pd_flag_stg0[0] || sc_flag_stg0[0]) && |PRD_rx_charisk[2:0]);
    // long starting in upper
    else if (PRD_idle2_selected && (pd_flag_stg0[1] || sc_flag_stg0[1]))
      control_sym_in_error_cond_dd[3] = |PRD_rx_charisk[6:1];
    // long starting in lower
    else if (PRD_idle2_selected && (pd_flag_stg0[0] || sc_flag_stg0[0] || lower_delimiter_q))
      control_sym_in_error_cond_dd[3] = ((lower_delimiter_q) && |PRD_rx_charisk[7:5]) ||
                                             ((pd_flag_stg0[0] || sc_flag_stg0[0]) && |PRD_rx_charisk[2:0]);
    else
      control_sym_in_error_cond_dd[3] = 1'b0;
  end

  // 4) Restart-from-Retry when not expecting one
  always @* begin
    if (rfr_detect_stg1)
      control_sym_in_error_cond_dd[4] = PR_input_status_good;
    else
      control_sym_in_error_cond_dd[4] = 1'b0;
  end

  // 5) Packet-Retry when in multi-VC mode
  // FIXVC
  //always @* begin                            // the control_sym_in_error_cond_dd[5] is always assigned to 0
  //  control_sym_in_error_cond_dd[5] = 1'b0;  // without left hand side operands, this loop is not activated
  //end                                        // To fix the CR 726266, this logic is commented and shifted in
                                               // 6) End-of-Packet when not in packet code part below

  //   6) End-of-Packet when not in packet
  always @* begin
    control_sym_in_error_cond_dd[6] = (|eop && ~|  in_packet_stg0) || &eop;
    control_sym_in_error_cond_dd[5] = 1'b0;    // To fix the CR 726266, this logic is added here
  end

  assign control_sym_in_error_cond_cmb = 
                                         |control_sym_in_error_cond_d;      // CR# 849355 fixed //

  assign control_sym_in_error_cond_dd_cmb = |control_sym_in_error_cond_dd;



  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      control_sym_in_error_cond_d   <= #TCQ 6'b0;
      prx_cs_in_error_cond          <= #TCQ 1'b0;
      control_sym_in_error_cond     <= #TCQ 1'b0;
      control_sym_in_error_straddle <= #TCQ 1'b0;
    end else begin
      control_sym_in_error_cond_d   <= #TCQ control_sym_in_error_cond_dd;
      prx_cs_in_error_cond          <= #TCQ |control_sym_in_error_cond_dd;
      control_sym_in_error_cond     <= #TCQ prx_cs_in_error_cond;
      control_sym_in_error_straddle <= #TCQ control_sym_in_error_straddle_d;
    end
  end

  // Specifically identify when there is a bad status symbol,
  // for use with link initializatin
  reg stat_q;
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      stat_q <= #TCQ 1'b0;
    end else begin
      stat_q <= #TCQ |stat;
    end
  end

  always @(posedge phy_clk) begin
    if (phy_rst_q)
      prx_rcvd_bad_status <= #TCQ 1'b0;
    else if (!pp_port_initialized_stg1 || PR_link_initialized)
      prx_rcvd_bad_status <= #TCQ 1'b0;
    else
      prx_rcvd_bad_status <= #TCQ (stat_q && |control_sym_in_error_cond_d[3:1]) || cs_crc_in_error_cond;
  end


  // In Retry Conditions -
  // 1) Receive a Stomp control symbol
  reg [1:0] lreq_q;
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      control_sym_retry_cond_d <= #TCQ 1'b0;
      control_sym_retry_cond   <= #TCQ 1'b0;
      lreq_q                   <= #TCQ 2'h0;
    end else begin
      control_sym_retry_cond_d <= #TCQ PR_input_status_good && |pd_flag_stg1 &&
                                       (stomp_detect_stg1 || (|(pd_flag_stg1 & lreq_q) && ~|lreq_in_stat_detect_stg1));
      control_sym_retry_cond   <= #TCQ control_sym_retry_cond_d;
      lreq_q                   <= #TCQ lreq;
    end
  end

 // for stomp, retry condition CR # 825747 is added
 wire control_sym_retry_cond_c;

 assign control_sym_retry_cond_c = PR_input_status_good && |pd_flag_stg1 &&
                                       (stomp_detect_stg1 || (|(pd_flag_stg1 & lreq_q) && ~|lreq_in_stat_detect_stg1));


    // *- COVERAGE (cp_PRX_long_cs_no_end_delimiter)
    // Observe a long control symbol with no end delimiter

    // *- COVERAGE (cp_PRX_long_cs_wrong_end_delimiter)
    // Observe a long control symbol with an end delimiter that doesn�t match the start delimiter

    // *- COVERAGE (cp_PRX_cs_bad_pd_delimiter)
    // Observe a PD start delimiter when SC should have been used

    // *- COVERAGE (cp_PRX_cs_bad_sc_delimiter)
    // Observe a SC start delimiter when PD should have been used

    // *- COVERAGE (cp_PRX_illegally_embedded_k_char)
    // Observe a control symbol with an illegally embedded K character

    // *- COVERAGE (cp_PRX_unexpected_rfr)
    // Observe a Restart-from-Retry when not in the Input Error stopped state

    // *- COVERAGE (cp_PRX_multi_vc_pr)
    // Observe a Packet-Retry when in multi-VC mode

    // *- COVERAGE (cp_PRX_non_consecutive_on_pa)
    // Observe a non-consecutive AckID on a Packet-Acknowledge

    // *- COVERAGE (cp_PRX_lresq_with_no_lreq)
    // Observe a Link-Response when no Link-Request was sent

    // *- COVERAGE (cp_PRX_non_consecutive_on_pr)
    // Observe a non-consecutive AckID on a Packet-Retry

    // *- COVERAGE (cp_PRX_non_consecutive_on_lresp)
    // Observe a non-consecutive AckID on a Link-Response (not an error)

    // *- COVERAGE (cp_PRX_unexpected_ackid_on_lresp)
    // Observe an unexpected AckID on a Link-Response (out_fatal)

    // *- COVERAGE (cp_PRX_lreq_coverage)
    // Observe a Link Request of type PD and SC in both IDLE1 and IDLE2

  // }}} End of Control Symbol Error ------


  // {{{ + IDLE Sequence Error Detection --
  // Checks being performed:
  // 1) Invalid IDLE1 sequence
  // 2) Invalid IDLE2 sequence
  integer ii;
  //wire [1:0] kchar_compare = {&PRD_rx_charisk[7:4], &PRD_rx_charisk[3:0]};
  reg  [7:0] idle1_compare, idle2_compare;
  reg  [1:0] idle_seq_in_error_cond_d;

  // only valid characters in IDLE1 = K, R, A
  // only valid characters in IDLE2 = K, R, A, M, and data
  always @* begin
    for (ii = 0; ii < 8; ii = ii + 1) begin
      idle1_compare[ii] = PRD_rx_data[ii*8 +: 8] == K_CHAR ||
                          PRD_rx_data[ii*8 +: 8] == R_CHAR ||
                          PRD_rx_data[ii*8 +: 8] == A_CHAR;
      idle2_compare[ii] = idle1_compare[ii] || PRD_rx_data[ii*8 +: 8] == M_CHAR;
    end
  end

  // only check IDLE patterns when not in a packet
  always @* begin
    if (PR_link_initialized) begin
      if (!in_packet_stg0[0] && !(pd_flag_stg0[0] || sc_flag_stg0[0])) begin
        if (PRD_idle2_selected && IDLE2)

          idle_seq_in_error_cond_d[0] = |(PRD_rx_charisk[3:0] & ~idle2_compare[3:0]) &&
                                        !(pd_flag_stg0[1] || sc_flag_stg0[1]);
        else // IDLE1
          idle_seq_in_error_cond_d[0] = !(&PRD_rx_charisk[3:0] && &idle1_compare[3:0]);
      end else begin
        idle_seq_in_error_cond_d[0] = 1'b0;
      end
      if (!in_packet_stg0[1] && !(pd_flag_stg0[1] || sc_flag_stg0[1])) begin
        if (PRD_idle2_selected && IDLE2)

          idle_seq_in_error_cond_d[1] = |(PRD_rx_charisk[7:4] & ~idle2_compare[7:4]) &&
                                        !(pd_flag_stg1[0] || sc_flag_stg1[0]);
        else // IDLE1
          idle_seq_in_error_cond_d[1] = !(&PRD_rx_charisk[7:4] && &idle1_compare[7:4]);
      end else begin
        idle_seq_in_error_cond_d[1] = 1'b0;
      end
    end else begin
      idle_seq_in_error_cond_d = 2'h0;
    end
  end

assign idle_seq_in_error_cond_cmb = idle_seq_in_error_cond_d; // 

  reg idle_seq_in_error_cond_stg1;//

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      idle_seq_in_error_cond_stg1 <= #TCQ 1'b0; // 
      idle_seq_in_error_cond      <= #TCQ 1'b0;
    end else begin
      idle_seq_in_error_cond_stg1 <= #TCQ |idle_seq_in_error_cond_d;// 
      idle_seq_in_error_cond      <= #TCQ idle_seq_in_error_cond_stg1;
    end
  end



    // *- COVERAGE (cp_PRX_idle1_char_error)
    // In IDLE1, observe an error on a K character,
    // while charisk is still asserted for that byte

    // *- COVERAGE (cp_PRX_idle1_m_error)
    // In IDLE1, observe an illegal /M/ character

    // *- COVERAGE (cp_PRX_idle1_no_charisk_error)
    // In IDLE1, observe a legally formed K character that does not have charisk asserted

    // *- COVERAGE (cp_PRX_idle2_char_error)
    // In IDLE2, observe an error on a K character,
    // while charisk is still asserted for that byte

    // *- COVERAGE (cp_PRX_idle2_no_charisk_error)
    // In IDLE2, observe a legally formed K character that does not have charisk asserted

  // }}} End of Idle Sequence Error -------

// detect invalid data characters in upper 32 bits of IDLE2, Part 6, section 5.13.2.2.2, 5.13.2.4
// // added to fix the CR # 842999
  wire [7:4] idle2_invalid_non_data_char_7_4;
  wire invalid_non_data_char_in_upper_32_bits;

  assign idle2_invalid_non_data_char_7_4[7] = PRD_rx_charisk[7] &&
                               (
                                (PRD_rx_data[63:56] == K_CHAR) // K_CHAR = BC
                                ||
                                (PRD_rx_data[63:56] == R_CHAR) // R_CHAR = FD
                                ||
                                (PRD_rx_data[63:56] == A_CHAR) // A_CHAR = FB
                               );

  assign idle2_invalid_non_data_char_7_4[6] = PRD_rx_charisk[6] &&
                               (
                                (PRD_rx_data[55:48] == K_CHAR) // K_CHAR = BC
                                ||
                                (PRD_rx_data[55:48] == R_CHAR) // R_CHAR = FD
                                ||
                                (PRD_rx_data[55:48] == A_CHAR) // A_CHAR = FB
                               );

  assign idle2_invalid_non_data_char_7_4[5] = PRD_rx_charisk[5] &&
                               (
                                (PRD_rx_data[47:40] == K_CHAR) // K_CHAR = BC
                                ||
                                (PRD_rx_data[47:40] == R_CHAR) // R_CHAR = FD
                                ||
                                (PRD_rx_data[47:40] == A_CHAR) // A_CHAR = FB
                               );

  assign idle2_invalid_non_data_char_7_4[4] = PRD_rx_charisk[4] &&
                               (
                                (PRD_rx_data[39:32] == K_CHAR) // K_CHAR = BC
                                ||
                                (PRD_rx_data[39:32] == R_CHAR) // R_CHAR = FD
                                ||
                                (PRD_rx_data[39:32] == A_CHAR) // A_CHAR = FB
                               );

  assign invalid_non_data_char_in_upper_32_bits = |idle2_invalid_non_data_char_7_4;

  // {{{ + Packet Error Detection ---------
  // Checks being performed:
  // 1) Packets that contain K characters, not part of embedded control symbols
  // 2) Packets that exceed the maximum packet length
  // 3) Packets whose CRC are not in the correct location
  reg  [3:1] packet_in_error_cond_d;

  // 1) Packets that contain K characters, not part of embedded control symbols
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      packet_in_error_cond_d[1] <= #TCQ 1'b0;
    end else if (!PR_link_initialized) begin
      packet_in_error_cond_d[1] <= #TCQ 1'b0;
    end else if (PRD_idle2_selected) begin
      if (in_packet_stg0[1]
          &&
          !(sc_flag_stg0[1] || pd_flag_stg0[1])
          &&
          !(sc_flag_stg1[0] || pd_flag_stg1[0])
          &&
          // this checks the upper 32 bit part of the data beats, if it has invlid characters
          invalid_non_data_char_in_upper_32_bits // added to fix the CR # 842999
          && // CR #820674, CR# 843008, Spec 6, sections 5.13.2.2.2, 5.13.2.4 //
             // added to fix idle2 based, if upper 32 bit part has errors, then it should be flagged even
          (idle2_sync_char_stg0 && |PRD_rx_charisk[3:0]) // though lower part starts with M (sync sequence)
          ) begin                                        // the above code checks the M in lower 32 data beats
        packet_in_error_cond_d[1] <= #TCQ 1'b1;
      end else if (in_packet_stg0[0]
                   &&
                   !(|sc_flag_stg0 || |pd_flag_stg0)
                   &&
                   |PRD_rx_charisk[3:0]  // this checks the lower 32 bit part of the data beats, CR# 843008, Spec 6, 5.13.2.2.2
                   &&                    // added to fix idle2 based
                   !idle2_sync_char_stg0 // CR #820674, as this is upper 32 bit part no need to check, the lower 32 bits
                   ) begin
        packet_in_error_cond_d[1] <= #TCQ 1'b1;
      end else begin
        packet_in_error_cond_d[1] <= #TCQ 1'b0;
      end
    end else begin
    if (packet_in_error_cond_d[1] == 1'b1) begin
        packet_in_error_cond_d[1] <= #TCQ 1'b0;
      end else if (in_packet_stg0[1] && !(sc_flag_stg0[1] || pd_flag_stg0[1]) && |PRD_rx_charisk[7:4]) begin
        packet_in_error_cond_d[1] <= #TCQ 1'b1;
      end else if (in_packet_stg0[0] && !(sc_flag_stg0[0] || pd_flag_stg0[0]) && |PRD_rx_charisk[3:0]) begin
        packet_in_error_cond_d[1] <= #TCQ 1'b1;
      end else begin
        packet_in_error_cond_d[1] <= #TCQ 1'b0;
      end
    end
  end


  // 2) Packets that exceed the maximum packet length -
  // The largest sized packet in this region is 276 bytes, which occupies 35 beats.
  reg [5:0] packet_length_count;
  always @* begin
    if (packet_length_count > 6'd35
            // added below condition while fixing CR #820674
            &&                    // The Sync Sequence in IDLE2, if its part of the packet followed by LREQ,
            !idle2_sync_char_stg1 // then the max packet length error should be supressed.
            )
      packet_in_error_cond_d[2] = 1'b1;
  else if ((packet_length_count == 6'd35)
            &&
            data_vld_stg1
            &&
            (!((ordered_rx_data_stg1[31:24] == (8'b01111100)) && lower_padded_stg1) | (PRD_idle2_selected && (carryover_stg2 ? data_vld_stg0_d[1] : data_vld_stg0_d[0])))
            &&
            (!((ordered_rx_data_stg1[31:24] == (8'b00011100)) && lower_padded_stg1) | (PRD_idle2_selected && (carryover_stg2 ? data_vld_stg0_d[1] : data_vld_stg0_d[0])))
            // added below condition while fixing CR #820674
            &&                    // The Sync Sequence in IDLE2, if its part of the packet followed by LREQ,
            !idle2_sync_char_stg1 // then the max packet length error should be supressed.
            )// CR 806709
      packet_in_error_cond_d[2] = 1'b1;
    else
      packet_in_error_cond_d[2] = 1'b0;
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q)
      packet_length_count <= #TCQ 6'h1;
    else if (PRD_idle2_selected && |(lreq) && |(in_packet_stg0)) // In IDLE2, if any LREQ is detected, at the end of packet
      packet_length_count <= #TCQ 6'h1;     // it means to cancell the packet.
    else if (framing_end_stg1)
      packet_length_count <= #TCQ 6'h1;
    else if (!PR_port_stat_ok)
      packet_length_count <= #TCQ 6'h1;
    else if (data_vld_stg1 && data_stream_enable_stg1)
      packet_length_count <= #TCQ packet_length_count + 1;
  end


  // 3) Packets whose CRC are not in the correct location
  // NOTE: This check was specifically added for cases where the expected location matches the crc check
  // but the actual CRC is elsewhere. This might be seen only in IDLE1, on b2b EOP, SOP where the
  // EOP is missing a charisk. This is very rare and will only need to be checked with the EOP and SOP
  // are reordered to show up on the same clock cycle of the ordered data.
  reg speculate_crc_loc_fail;
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      speculate_crc_loc_fail <= #TCQ 1'b0;
    end else if (data_vld_stg1) begin
      speculate_crc_loc_fail <= #TCQ |crc_loc_stg1[3:2] && !lower_padded_stg1;
    end
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      packet_in_error_cond_d[3] <= #TCQ 1'b0;
    end else if (!PR_link_initialized) begin
      packet_in_error_cond_d[3] <= #TCQ 1'b0;
    end else begin
      if (framing_end_stg1 && !framing_dsc_stg1 && data_vld_stg1 && !first_beat_stg1 &&
          rt_stream_enable_stg2 && |crc_loc_stg1[3:2] && !lower_padded_stg1) begin
        packet_in_error_cond_d[3] <= #TCQ 1'b1;
      end else if (framing_end_stg1 && !framing_dsc_stg1 && !data_vld_stg1 &&
                   rt_stream_enable_stg2 && |crc_loc_stg1[3:2]) begin
        packet_in_error_cond_d[3] <= #TCQ speculate_crc_loc_fail;
      end else begin
        packet_in_error_cond_d[3] <= #TCQ 1'b0;
      end
    end
  end


  always @(posedge phy_clk) begin
    if (phy_rst_q)
      packet_in_error_cond <= #TCQ 1'b0;
    else
      packet_in_error_cond <= #TCQ |packet_in_error_cond_d;
  end

    // *- COVERAGE (cp_PRX_k_char_in_packet)
    // Observe a K character in the middle of a packet, that is not part of an embedded control symbol

    // *- COVERAGE (cp_PRX_packet_too_long)
    // Observe a packet whose length exceeds the maximum

  // }}} End of Packet Error Detection ----


  // {{{ + CRC Check ----------------------
  // Checks being performed:
  // 1) Control symbol with a bad CRC
  // 2) Packet with a bad mid-CRC
  // 3) packet with a bad final CRC


  // 1) Control symbol with a bad CRC

  // short upper
  wire [18:0] short_cs_fields_0     = PRD_rx_data[55:37];
  wire  [4:0] short_cs_actual_crc_0 = PRD_rx_data[36:32];
  wire  [4:0] short_cs_expected_crc_0;
  srio_gen2_v4_1_16_crc5_20 short_crc_cs0_inst
    (.crc    (short_cs_expected_crc_0),
     .din    (short_cs_fields_0));

  // short lower
  wire [18:0] short_cs_fields_1     = PRD_rx_data[23:5];
  wire  [4:0] short_cs_actual_crc_1 = PRD_rx_data[4:0];
  wire  [4:0] short_cs_expected_crc_1;
  srio_gen2_v4_1_16_crc5_20 short_crc_cs1_inst
    (.crc    (short_cs_expected_crc_1),
     .din    (short_cs_fields_1));

  // long upper
  wire [34:0] long_cs_fields_0     = PRD_rx_data[55:21];
  wire [12:0] long_cs_actual_crc_0 = PRD_rx_data[20:8];
  wire [12:0] long_cs_expected_crc_0;
  srio_gen2_v4_1_16_crc13_35 long_crc_cs0_inst
    (.crc    (long_cs_expected_crc_0),
     .din    (long_cs_fields_0));
  // long lower
  wire [23:0] long_cs_first_half_1 = PRD_rx_data[23:0];
  reg  [23:0] long_cs_first_half_1_q;
  always @(posedge phy_clk) begin
    long_cs_first_half_1_q <= #TCQ long_cs_first_half_1;
  end

  wire [34:0] long_cs_fields_1     = {long_cs_first_half_1_q, PRD_rx_data[63:53]};
  wire [12:0] long_cs_actual_crc_1 = PRD_rx_data[52:40];
  wire [12:0] long_cs_expected_crc_1;
  srio_gen2_v4_1_16_crc13_35 long_crc_cs1_inst
    (.crc    (long_cs_expected_crc_1),
     .din    (long_cs_fields_1));

  always @(posedge phy_clk) begin
    cs_crc_in_error_cond         <= #TCQ |prx_cs_crc_check_fail;
    cs_crc_in_error_cond_mod     <= #TCQ |prx_cs_crc_check_fail[2:0];
    cs_crc_in_error_cond_mod_q   <= #TCQ cs_crc_in_error_cond_mod;

    // crc error in upper, IDLE1
    prx_cs_crc_check_fail[0]     <= #TCQ (pd_flag_stg0[1] || sc_flag_stg0[1]) && !PRD_idle2_selected &&
                                         (short_cs_expected_crc_0 != short_cs_actual_crc_0);
    // crc error in lower, IDLE1
    // special case for when there is an eop and sop in the same beat, where the sop has an error.
    // Delay the detection of this scenario by one cycle to avoid interfering with the previous packet.
    prx_cs_crc_check_fail[1]     <= #TCQ ((pd_flag_stg0[0] || sc_flag_stg0[0]) && !PRD_idle2_selected &&
                                         (short_cs_expected_crc_1 != short_cs_actual_crc_1) && !(eop[1] && sop[0])) ||
                                         prx_cs_crc_check_fail_early;
    prx_cs_crc_check_fail_early  <= #TCQ ((pd_flag_stg0[0] || sc_flag_stg0[0]) && !PRD_idle2_selected &&
                                         (short_cs_expected_crc_1 != short_cs_actual_crc_1) && (eop[1] && sop[0]));
    // crc error in upper, IDLE2
    prx_cs_crc_check_fail[2]     <= #TCQ (pd_flag_stg0[1] || sc_flag_stg0[1]) && PRD_idle2_selected &&
                                         (long_cs_expected_crc_0 != long_cs_actual_crc_0);
    // crc error in lower, IDLE2
    prx_cs_crc_check_fail[3]     <= #TCQ (pd_flag_stg1[0] || sc_flag_stg1[0]) && PRD_idle2_selected &&
                                         (long_cs_expected_crc_1 != long_cs_actual_crc_1);
    prx_cs_crc_check_fail_q      <= #TCQ prx_cs_crc_check_fail;
  end

  // 2) Packet with a bad mid-CRC
  // 3) packet with a bad final CRC

  // Generate the CRC value for the incoming packet. No reset is needed
  // because it resets on every SOF before use.
  wire  [15:0] crc16_d, crc32_d, crc48_d, crc64_d;
  reg   [15:0] crc64;

  // Register the outputs
  // Calculate the value of the CRC for various valid bytes
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      crc64 <= #TCQ 16'hFFFF;
    end else if (framing_end_stg1 || !PR_port_stat_ok) begin
      crc64 <= #TCQ 16'hFFFF;
    end else if (data_vld_stg1) begin
      crc64 <= #TCQ crc64_d;
    end
  end

  // 16-bit wide Next CRC Combinational Equations
  srio_gen2_v4_1_16_crc16_16 ollm_rx_crc16_16_inst (
    .din   (masked_rx_data_stg1[63:48]),
    .cin   (crc64),
    .crc   (crc16_d)
  );

  // 32-bit wide Next CRC Combinational Equations
  srio_gen2_v4_1_16_crc16_32 ollm_rx_crc16_32_inst (
    .din   (masked_rx_data_stg1[63:32]),
    .cin   (crc64),
    .crc   (crc32_d)
  );

  // 48-bit wide Next CRC Combinational Equations
  srio_gen2_v4_1_16_crc16_48 ollm_rx_crc16_48_inst (
    .din   (masked_rx_data_stg1[63:16]),
    .cin   (crc64),
    .crc   (crc48_d)
  );

  // 64-bit wide Next CRC Combinational Equations
  srio_gen2_v4_1_16_crc16_64 ollm_rx_crc16_64_inst (
    .din   (masked_rx_data_stg1),
    .cin   (crc64),
    .crc   (crc64_d)
  );


  // registered earlier to improve timing. So, this is combinatorial.
  reg       pk_crc_in_error_cond_d;
  reg       pk_crc_in_error_cond_standard_case;
  reg       pk_crc_in_error_cond_standard_condition;
  reg [8:1] pk_crc_in_error_cond_speculate;
  reg       single_cycle_pkt;
  always @* begin
    case (crc_loc_stg1)
    4'b1000 : pk_crc_in_error_cond_d = (crc64 != masked_rx_data_stg1[63:48]);
    4'b0100 : pk_crc_in_error_cond_d = (crc16_d != masked_rx_data_stg1[47:32]);
    4'b0010 : pk_crc_in_error_cond_d = (crc32_d != masked_rx_data_stg1[31:16]);

    default : pk_crc_in_error_cond_d = (crc48_d != masked_rx_data_stg1[15:0]);

    endcase
  end
  always @(posedge phy_clk) begin
    pk_crc_in_error_cond_standard_case <= #TCQ pk_crc_in_error_cond_d;
    pk_crc_in_error_cond_standard_condition <= #TCQ framing_end_stg1 && data_vld_stg1 && !first_beat_stg1
                                                    ;
  end
  always @(posedge phy_clk) begin
    if(PRD_idle2_selected && (idle2_sync_char_stg0 && |PRD_rx_charisk[3:0]))       // updated to (idle2_sync_char_stg0 && |PRD_rx_charisk[3:0])
      pk_crc_in_error_cond_speculate    <= 7'b0;         //                           the above chage allows to detect errors in upper 32 bits of data beat
    else if (data_vld_stg1) begin
      pk_crc_in_error_cond_speculate[8] <= #TCQ (crc64 != masked_rx_data_stg1[63:48]);
      pk_crc_in_error_cond_speculate[4] <= #TCQ (crc16_d != masked_rx_data_stg1[47:32]);
      pk_crc_in_error_cond_speculate[2] <= #TCQ (crc32_d != masked_rx_data_stg1[31:16]);
      pk_crc_in_error_cond_speculate[1] <= #TCQ (crc48_d != masked_rx_data_stg1[15:0]);
    end
  end

  // single-cycle packets have to be treated a bit differently because
  // the crc location hasn't been determined yet.
  always @(posedge phy_clk) begin
    if (phy_rst_q)
      single_cycle_pkt <= #TCQ 1'b0;
    else
      single_cycle_pkt <= #TCQ framing_end_stg1 && data_vld_stg1 && first_beat_stg1;
  end

wire crc_check; // Fix for CR# 847695
wire  [15:0] crc48_check;
  // 16-bit wide Next CRC Combinational Equations
  srio_gen2_v4_1_16_crc16_48 ollm_rx_crc48_check_inst (
    .din   (masked_rx_data_stg1[63:16]),
    .cin   (crc64),
    .crc   (crc48_check)
  );

wire  [15:0] crc32_check;
  // 16-bit wide Next CRC Combinational Equations
  srio_gen2_v4_1_16_crc16_32 ollm_rx_crc16_check_inst (
    .din   (masked_rx_data_stg1[63:32]),
    .cin   (crc64),
    .crc   (crc32_check)
  );


reg [1:0] sop_reg;
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      sop_reg <= #TCQ 2'b0;
    end else begin
      sop_reg <= #TCQ sop;
    end
  end

wire crc_issue_48_bit;
assign crc_issue_48_bit = (crc48_check != masked_rx_data_stg1[15:0])? 1'b1:1'b0;

wire crc_issue_32_bit;
assign crc_issue_32_bit = (crc32_check != masked_rx_data_stg1[31:16])? 1'b1:1'b0;

wire masked_data_padded_with_0;
assign masked_data_padded_with_0 = !(|masked_rx_data_stg1[15:0])? 1'b0:1'b1;

wire catch_crc_error;
assign catch_crc_error = !(|masked_rx_data_stg1[15:0])? crc_issue_32_bit : crc_issue_48_bit;

assign crc_check = (PRD_idle2_selected 
                    && 
		    PR_link_initialized 
		    && 

		    catch_crc_error
		    && 
		    pd_flag_stg1[0]
		    &&
		    PRD_rx_charisk_reg2[4]
		    &&
		    PRD_rx_charisk_reg[3]
		    &&
		    |in_packet_stg0
		    &&
		    data_vld_stg1//
		    &&
		    //
		    framing_end_stg1
		    &&
		    sop_reg[0]
		    &&
            idle2_sync_char_stg0
		    &&
		    masked_data_padded_with_0
		    )?
		   1'b1:
		   1'b0;

reg crc_check_reg;
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      crc_check_reg <= #TCQ 1'b0;
    end else begin
      crc_check_reg <= #TCQ crc_check;
    end
  end

  reg pk_crc_in_error_cond_raw;
  assign pk_crc_in_error_cond = (PRD_idle2_selected && idle2_sync_char_stg2)?// updated from idle2_sync_char_stg0 to idle2_sync_char_stg2 to fix CR# 847208 and CR# 847695, //
                                 1'b0                                         // this is combo logic and will restrict only to stg2 use only for the current packet 
                                 :
                                (
                                  pk_crc_in_error_cond_standard_condition?
                                  ( pk_crc_in_error_cond_standard_case  | 
  				                   (pk_crc_in_error_cond_raw && data_stream_enable_stg1)
				                   )
                                   :
                                  (pk_crc_in_error_cond_raw && data_stream_enable_stg1)
				 ||
				 crc_check_reg // Fix for CR# 847695
                                );

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      pk_crc_in_error_cond_raw <= #TCQ 1'b0;
    // below "idle2_sync_char_stg0" condition is applicable only for IDLE2 cases //
    // when IDLE2 sync sequence is detected, LREQ would be followed
    // the packet should be considered as cancelled and no errors should be reported
    // as per discussion with Barry Richard, core should not generate any error and enter into Retry Stopped State
    // Page 153, Spec 6 - "The cancellation of a packet shall not result in the generation or report of any errors."
    //end else if (idle2_sync_char_stg0 || |(lreq)) begin // 
    //end else if (idle2_sync_char_stg0 || |(lreq)) begin // 
    end else if (PRD_idle2_selected && |(lreq)) begin // 
      pk_crc_in_error_cond_raw <= #TCQ 1'b0; // 
    // if framing_end shows up some number of cycles after the last valid data
    end else if (framing_end_stg1 && !data_vld_stg1 && beat_count_q_is_10 && !mid_crc_loc_stg1) begin
      pk_crc_in_error_cond_raw <= #TCQ pk_crc_in_error_cond_speculate[crc_loc_stg2];
    // if it's a single cycle or if the last beat comes without data
    end else if (!ignore_pk_crc && ((single_cycle_pkt && !framing_dsc_stg1_delay)|| (framing_end_stg1 && !data_vld_stg1))) begin
      pk_crc_in_error_cond_raw <= #TCQ pk_crc_in_error_cond_speculate[crc_loc_stg1];
    // confirm that the mid_crc is correct
    end else if (mid_crc_loc_stg1 && !mid_crc_loc_stg2) begin
      pk_crc_in_error_cond_raw <= #TCQ (crc64 != masked_rx_data_stg1[63:48])
                                       &&
                                      !(PRD_idle2_selected && // 
                                        (idle2_sync_char_stg0 && |PRD_rx_charisk[3:0]));// updated to make sure to detect all upper
                                                                                        // 32 bit data beat errors

    end else begin
      pk_crc_in_error_cond_raw <= #TCQ 1'b0;
    end
  end

/*  reg [1:0] sop_stg1;
    reg [1:0] eop_stg1;
*/
  reg sop_stg1;
  reg eop_stg1;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      sop_stg1   <= #TCQ 1'b0;
      eop_stg1   <= #TCQ 1'b0;
  /*  sop_stg1   <= #TCQ 2'b0;
      eop_stg1   <= #TCQ 2'b0;
  */
      framing_dsc_stg1_delay   <= #TCQ 1'b0;
    end else begin
      sop_stg1   <= #TCQ |sop;
      eop_stg1   <= #TCQ |eop;
      /*sop_stg1   <= #TCQ sop;
      eop_stg1   <= #TCQ eop;
      */
      framing_dsc_stg1_delay   <= #TCQ framing_dsc_stg1;
    end
  end

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      ignore_pk_crc   <= #TCQ 1'b0;
    end else begin
      ignore_pk_crc   <= #TCQ prx_in_retry_detect || control_sym_retry_cond_c || control_sym_retry_cond_d || // added || control_sym_retry_cond_c, CR# 825747
                              (
                              (stomp_detect_stg1
                              || (lreq_detect_stg1 && !eop_stg1 && !sop_stg1)       // 
                              )
                              && !single_cycle_pkt
                              );
    end
  end

  assign crc_in_error_cond = cs_crc_in_error_cond_mod_q || (pk_crc_in_error_cond && !ignore_pk_crc && PR_port_stat_ok);


    // *- COVERAGE (cp_PRX_bad_mid_crc)
    // Observe a bad mid-term packet CRC

    // *- COVERAGE (cp_PRX_bad_final_crc)
    // Observe a bad final packet CRC

    // *- COVERAGE (cp_PRX_bad_short_cs_crc)
    // Observe a bad short control symbol CRC

    // *- COVERAGE (cp_PRX_bad_long_cs_crc)
    // Observe a bad long control symbol CRC

  // }}} End of CRC Check -----------------
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
        rx_charisk_stg1 <= 4'b0;
    end else begin
        rx_charisk_stg1 <= {PRD_rx_charisk[7],
                            PRD_rx_charisk[4],
                            PRD_rx_charisk[3],
                            PRD_rx_charisk[0]} ;
    end
  end


  // {{{ + AckID Check --------------------
  // Checks being performed:
  // 1) Packet with unexpected AckID (must increment by one every time)
  wire [5:0] received_ackid;
  generate if (IDLE2 == 1) begin : received_ackid_idle2_gen
    assign received_ackid = PRD_idle2_selected ? ordered_rx_data_stg1[63:58]
                            : {1'b0, ordered_rx_data_stg1[63:59]};
  end else  begin                : received_ackid_idle1_gen
    assign received_ackid[5:0] = {1'b0, ordered_rx_data_stg1[63:59]};
  end
  endgenerate
  wire [5:0] prx_next_rcvd_pkt_int;
  reg  [5:0] prx_next_rcvd_pkt_int_full;
  reg  [5:0] prx_next_rcvd_pkt_full, prx_last_good_pkt_full;

  // update the next expected AckID value once the packet exits without any errors detected
  // for every framing end we see with no prevailing errors or retries, increment
  // the next expected value and the last good packet value for the OLLM TX
  assign PRX_next_rcvd_pkt     = {PRD_idle2_selected && prx_next_rcvd_pkt_full[5], prx_next_rcvd_pkt_full[4:0]};
  assign prx_next_rcvd_pkt_int = {PRD_idle2_selected && prx_next_rcvd_pkt_int_full[5], prx_next_rcvd_pkt_int_full[4:0]};
  assign PRX_last_good_pkt     = {PRD_idle2_selected && prx_last_good_pkt_full[5], prx_last_good_pkt_full[4:0]};
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      prx_next_rcvd_pkt_full     <= #TCQ 6'h00;
      prx_next_rcvd_pkt_int_full <= #TCQ 6'h00;
      prx_last_good_pkt_full     <= #TCQ 6'h3F;
    end else if (PC_load_nextpkt) begin
      prx_next_rcvd_pkt_full     <= #TCQ PC_next_rcvd_pkt;
      prx_next_rcvd_pkt_int_full <= #TCQ PC_next_rcvd_pkt;
      prx_last_good_pkt_full     <= #TCQ PC_next_rcvd_pkt - 1;
    end else begin
      if (framing_end_stg1      &&
                   rt_stream_enable_stg2 &&
                   !prx_in_retry_detect  &&
                   !prx_in_recoverable_detect &&
                   !framing_dsc_stg1     &&
                   !(first_valid_beat_stg1 && (rx_buf_retry_cond_d || control_sym_retry_cond_d))
                   ) begin
        prx_next_rcvd_pkt_int_full <= #TCQ prx_next_rcvd_pkt_int_full + 1;
      end else if (!PR_port_stat_ok
                  || prx_in_recoverable_detect // CR# 822485, in any recoverable error case, revert to next expected pkt_id
                  ) begin
        prx_next_rcvd_pkt_int_full <= #TCQ prx_next_rcvd_pkt_full;
      end
      if (PR_phyr_tvalid && BR_phyr_tready && PR_phyr_tlast && !PR_phyr_tuser[0]) begin
        if (PRD_idle2_selected) begin
          prx_last_good_pkt_full      <= #TCQ prx_last_good_pkt_full + 1;
          prx_next_rcvd_pkt_full      <= #TCQ prx_next_rcvd_pkt_full + 1;
        end else begin
          prx_last_good_pkt_full[4:0] <= #TCQ prx_last_good_pkt_full + 1;
          prx_last_good_pkt_full[5]   <= #TCQ 1'b0;
          prx_next_rcvd_pkt_full[4:0] <= #TCQ prx_next_rcvd_pkt_full + 1;
          prx_next_rcvd_pkt_full[5]   <= #TCQ 1'b0;
        end
      end
    end
  end


  // final determination if there is an error in the expected AckID
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      ackid_in_error_cond <= #TCQ 1'b0;
    end else if (first_valid_beat_stg1
                 &&
                 PR_port_stat_ok
                 &&
                 !(prx_in_retry_detect
                   ||
                   prx_in_retry_detect_q
                   ||
                   control_sym_retry_cond_d
                   )
                 &&                   // added to fix idle2 based
                 !idle2_sync_char_stg1// CR #820674
                 &&                                                // added to fix the CR 837145, when LREQ+RST/STATUS is
                 !(PRD_idle2_selected && |(lreq)) // present, dont detect the ackid errors
                 ) begin
      if (prx_next_rcvd_pkt_int != received_ackid) begin
        ackid_in_error_cond <= #TCQ 1'b1;
      end else begin
        ackid_in_error_cond <= #TCQ 1'b0;
      end
    end else begin
      ackid_in_error_cond <= #TCQ 1'b0;
    end
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      ackid_in_error_cond_q <= #TCQ 1'b0;
    end else begin
      ackid_in_error_cond_q <= #TCQ ackid_in_error_cond;
    end
  end


    // *- COVERAGE (cp_PRX_unexpected_ackid)
    // Observe an incoming packet with an unexpected AckID

    // *- COVERAGE (cp_PRX_last_good_pkt_during_error)
    // Observe the conditions under which last_good_pkt increments at the same time
    // as an error or retry condition

    // *- COVERAGE (cp_PRX_last_good_pkt_1after_error)
    // Observe the conditions under which last_good_pkt increments one cycle after
    // an error or retry condition

    // *- COVERAGE (cp_PRX_last_good_pkt_1before_error)
    // Observe the conditions under which last_good_pkt increments one cycle before
    // an error or retry condition

  // }}} End of AckID Check ---------------


  // {{{ + RX Buf Overflow Prevention -----
  // Checks being performed:
  // 1) Does the buffer have enough space for a packet of a given priority?
  // 2) RX Buffer drops TREADY, causing a source discontinue
  wire [1:0] packet_priority = ordered_rx_data_stg1[55:54];
  wire       response_type = ordered_rx_data_stg1[51:48] == 4'd13;

  assign rx_buf_retry_cond_d = BR_phy_buf_stat == 6'h00 ? 1'b1 :
                               BR_phy_buf_stat == 6'h01 ? (packet_priority < 2'h3) || (response_type != 1) :
                               BR_phy_buf_stat == 6'h02 ? packet_priority < 2'h2 :
                               BR_phy_buf_stat == 6'h03 ? packet_priority < 2'h1 :
                                                          1'b0;

  reg pr_port_retry;
  always @(posedge phy_clk) begin
    pr_port_retry <= #TCQ PR_port_stat == PORT_STAT_RETRY_STOP;
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q)
      rx_buf_retry_cond <= #TCQ 1'b0;
    else if (!pp_port_initialized_stg1)
      rx_buf_retry_cond <= #TCQ 1'b0;
    else if (dest_dsc_stg2 && !pr_port_retry)
      rx_buf_retry_cond <= #TCQ 1'b1;
    else if (first_valid_beat_stg1)
      rx_buf_retry_cond <= #TCQ rx_buf_retry_cond_d;
    else
      rx_buf_retry_cond <= #TCQ 1'b0;
  end


    // *- COVERAGE (cp_PRX_buf_stat_cross_priority)
    // Cross all priorities crossed with buf_stat {0, 1, 2, 3, 4+},
    // crossed with all VCs

  // }}} End of RX Buf Overflow -----------


  // {{{ + Other Error Detection ----------
  // Checks being performed:
  // 1) In maintenance-only mode, receive a non-maintenance packet
  // 2) Scrambler out of sync (from OPLM)
  reg  [2:1] other_in_error_cond_d;


  // 1) In maintenance-only mode, receive a non-maintenance packet
  always @* begin
    if (PC_input_maint_only && (first_valid_beat_stg1))
      other_in_error_cond_d[1] = ordered_rx_data_stg1[51:48] != FTYPE_MAINT;
    else
      other_in_error_cond_d[1] = 1'b0;
  end

  // 2) Scrambler out of sync (from OPLM)
  always @* begin
    if (pp_port_initialized_stg1 && pp_out_of_sync_stg1)
      other_in_error_cond_d[2] = 1'b1;
    else
      other_in_error_cond_d[2] = 1'b0;
  end

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      other_in_error_cond   <= #TCQ 1'b0;
      loss_of_sync          <= #TCQ 1'b0;
      rcvd_non_maint_packet <= #TCQ 1'b0;
    end else begin
      other_in_error_cond   <= #TCQ |other_in_error_cond_d;
      loss_of_sync          <= #TCQ other_in_error_cond_d[2];
      rcvd_non_maint_packet <= #TCQ other_in_error_cond_d[1];
    end
  end


    // *- COVERAGE (cp_PRX_unexpected_non_maint)
    // Observe a non-maintenance packet when in maintenance-only mode

    // *- COVERAGE (cp_PRX_expected_maint)
    // Observe a maintenance packet when in maintenance-only mode

    // *- COVERAGE (cp_PRX_out_of_sync)
    // Observe an out of sync error


  // }}} End of Other Error Detection -----

  // }}} End classes of error detections --

endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
//
// OLLM_RX_TOP
// Description:
// This module instantiates all the submodules of the OLLM RX design
//
// Hierarchy:
// PHY_TOP
//    |___OLLM_RX_TOP <-- this module
//             |_____OLLM_RX_CS_DECODE
//             |_____OLLM_RX_DATAPATH
//             |_____OLLM_RX_ERR_DETECT
// ---------------------------------------------------------------------

`timescale 1ps/1ps

module srio_gen2_v4_1_16_ollm_rx_top
  #(
    parameter TCQ           = 100,  // in pS
    parameter IDLE1         = 1,    // Include the IDLE1 sequence {0, 1}
    parameter IDLE2         = 0,    // Include the IDLE2 sequence {0, 1}
    parameter MODE_XG       = 5,    // Line rates {1/1.25, 2/2.5, 3/3.125, 5/5, 6/6.25}
    parameter VC            = 0,    // Highest number VC supported {0, 1}
    parameter SWITCH_MODE   = 0,    // If the core is generated with Switch Mode Support {0, 1}
    parameter RETRY         = 1,    // Includes Retry protocol {0, 1}
    parameter TARGET_DS     = 0, 
    parameter LINK_REQUESTS = 3,    // Additional link requests to send prior to port_error {0, 1, 2, 3, 4, 5, 6, 7}
    parameter VC1_CT        = 1,    // Default traffic mode for VC1 {0, 1}
    parameter LINK_WIDTH    = 1)
   (
  // {{{ port declarations ----------------
    // clocks and resets and general signals
    input             phy_clk,                    // PHY interface clock
    input             phy_rst,                    // Reset for PHY clock Domain
    input             log_clk,                    // LOG interface clock
    input             log_rst,                    // Reset for LOG clock Domain
    input             gt_pcs_clk,                 // GT interface clock
    output            PR_phy_rcvd_mce,            // MCE control symbol received
    output            PR_phy_rcvd_link_reset,     // Received 4 consecutive link reset control symbols
    output     [63:0] PR_debug,                   // OLLM RX Debug bus, should include useful signals for HW debug

    // OPLM Interface
    input      [63:0] PP_rx_data,                 // Receive data
    input      [7:0]  PP_rx_charisk,              // Indicates which bytes are K characters
    input      [1:0]  PP_rx_valid,                // Indicates valid words
    input             PP_idle2_selected,          // Indicates when an IDLE2 sequence is present
    input             PP_out_of_sync,             // Scrambler is out of sync
    input             PP_port_initialized,        // Indicates port is initialized
    input             PP_mode_1x,                 // Indicates the link trained down to 1x
    input      [LINK_WIDTH*4-1:0] PP_gt_decode_error,   // INVALID on GT RX (notintable or disperr)


    // RX Buffer Interface
    output            PR_phyr_tvalid,             // Valid data indicator
    input             BR_phyr_tready,             // Destination Ready
    output     [63:0] PR_phyr_tdata,              // Packet for transfer
    output     [7:0]  PR_phyr_tkeep,              // Byte Enable for transferred packet
    output            PR_phyr_tlast,              // Last DW of incoming packet
    output     [7:0]  PR_phyr_tuser,              // {1'b0, skip_crc, 3'h0, VC, CRF, src_dsc} AXI Compliance Pad
    input      [5:0]  BR_phy_buf_stat,            // Buffer status from the RX Buffer

    // OLLM TX Interface
    input             PT_sent_init_cs,            // Indicates we sent 15 control symbols
    output            PR_link_initialized,        // Indicates we are ready to transmit data
    output            PR_rewind,                  // An error or retry condition has been seen
    output     [5:0]  PR_phy_last_ack,            // Last PA received by the PHY core
    input      [5:0]  PT_phy_next_fm,             // Next Packet's Ack ID
    output     [5:0]  PR_phy_rcvd_buf_stat,       // Buffer status received from the link partner
    output            PR_send_rfr,                // Send an RFR control symbol (Request)
    input             PT_rfr_sent,                // Sent RFR (Grant)
    output            PR_send_lreq,               // Send a Link Request Control Symbol
    input             PT_lreq_sent,               // Sent Link Request
    output            PR_send_pna,                // Send a PNA control symbol
    input             PT_pna_sent,                // Sent PNA
    output            PR_send_pr,                 // Send a PR control symbol
    input             PT_pr_sent,                 // Sent PR
    output            PR_send_lresp,              // Send a Link Response Control Symbol
    input             PT_lresp_sent,              // Sent Link Response
    output     [4:0]  PR_cause,                   // Last cause for a PNA to send
    output     [4:0]  PR_port_stat,               // Current port status
    output     [5:0]  PR_last_good_pkt,           // Last PA to send
    output            PR_output_retry_stop,       // OLLM RX is currently in Output Retry Stopped State
    output            PR_output_error_stop,       // OLLM RX is currently in Output Error Stopped State
    output            PR_port_error,              // OLLM RX is currently in Port Error State
    output            PR_input_retry_stop,        // OLLM RX is currently in Input Retry Stopped State
    output            PR_input_error_stop,        // OLLM RX is currently in Input Error Stopped State
    output            PR_rcvd_error_free_status,  // Asserts when an error free status control symbol is received
    input             PT_sample_next_fm,          // Indicates to the ollm rx to sample the next fm

    // PHY Config Interface
    input      [5:0]  PC_next_rcvd_pkt,           // Load value for Next Expected packet
    input      [5:0]  PC_last_ack,                // Load value for phy_last_ack when Pload_ackids is asserted
    input             PC_load_ackids,             // Loads next_rcvd_pkt and last_ack with the CFG provided alternatives
    input             PC_load_nextpkt,            // Load next_rcvd_pkt with CFG value
    input             PC_send_lreq,               // Send a Link Request Input Status CS
    input       [2:0] PC_lreq_cmd,                // Command information for PC_send_lreq
    input      [23:0] PC_link_timeout,            // Time-out value for packet acknowledgement
    input             PC_clr_port_error,          // Clear the Output port error state
    input             PC_input_maint_only,        // Only maintenance traffic is allowed
    input             PC_error_disable,           // Disable error checking in the OLLM RX
// FIXVC - next two signals currently unused
    input             PC_vc_ct,                   // VC1 is in continuous traffic mode and all VC1 should be acked
    input             PC_vc_en,                   // Enable VC1 operation
    output            PR_rcvd_lresp,              // Asserted when a link response has been received
    output     [5:0]  PR_ackid_status,            // ackid status field from an LRESP
    output     [4:0]  PR_rcvd_port_stat,          // Last received link partner's port status
    output     [5:0]  PR_next_rcvd_pkt,           // Next expected packet AckID
    output            PR_rcvd_pa_or_pna           // Asserted when a Packet Accepted or Not Accepted has been received
  // }}} ----------------------------------
   );

  // {{{ wire declarations ----------------
  // Prefix notation:
  // phy = phy clock domain
  // pr/PR = Physical Layer Receive
  // pt/PT = Physical Layer Transmit
  // pc/PC = Physical Layer Config
  // pp/PP = Physical Layer OPLM
  // br/BR = Buffer Layer Receive
  // prx   = Physical Layer Error Detection signals (Not 'pre' to avoid confusion)
  // _st*  = Pipeline Stage Number

  // resets
  reg                    phy_rst_q = 1;              // registered physical layer reset
  reg                    log_rst_q = 1;              // registered logical layer reset

  // OLLM Decode Interface
  wire  [63:0]           prd_rx_data;                // Receive data
  wire  [7:0]            prd_rx_charisk;             // Indicates which bytes are K characters
  wire  [1:0]            prd_rx_valid;               // Indicates valid words
  wire                   prd_idle2_selected;         // Indicates when an IDLE2 sequence is present
  wire  [81:0]           prd_cs_decode;              // A whole series of control symbol decodes. See assignment

  // Pipeline stage 0 signals
  // - Data Parser
  wire  [1:0]            pd_flag_stg0;               // Packet Delimiter Delimiter indication
  wire  [1:0]            sc_flag_stg0;               // Control Symbol Delimiter indication

  // - Stype1 Decode
  wire  [1:0]            in_packet_stg0;             // indicates when the the data stream is part of a packet
  wire  [1:0]            sop;                        // successful decode of SOP in either upper or lower
  wire  [1:0]            stomp;                      // successful decode of STOMP in either upper or lower
  wire  [1:0]            eop;                        // successful decode of EOP in either upper or lower
  wire  [1:0]            rfr;                        // successful decode of RFR in either upper or lower
  wire  [1:0]            lreq;                       // successful decode of LREQ in either upper or lower
  wire  [1:0]            mce;                        // successful decode of MCE in either upper or lower

  // - Stype0 Decode
  wire  [1:0]            stat;                       // successful decode of STATUS in either upper or lower


  // Pipeline stage 1 signals
  // - Carryover from Stage 0
  wire                   pp_out_of_sync_stg1;        // Scrambler is out of sync
  wire                   pp_port_initialized_stg1;   // Indicates port is initialized

  wire                   framing_start_stg1;         // used with in_packet to indicate the start of a packet
  wire                   framing_end_stg1;           // used with in_packet to indicate the end of a packet
  wire                   framing_dsc_stg1;           // used with in_packet to indicate a discontinued packet
  wire  [5:0]            pa_ackid_stg1;              // sampled from parameter0 - pa ackid
  wire  [5:0]            pr_ackid_stg1;              // sampled from parameter0 - pr ackid
  wire                   lreq_detect_stg1;           // Link-Request detection
  wire  [1:0]            lreq_in_stat_detect_stg1;   // Link-Request detection - in stat
  wire                   lresp_detect_stg2;          // Link-Response detection
  wire                   rfr_detect_stg1;            // RFR detection
  wire                   pr_detect_stg1;             // PR detection
  wire  [1:0]            pa_detect_stg1;             // PA detection
  wire                   stomp_detect_stg1;          // PA detection
  wire  [1:0]            expected_ackid_coef_stg1;   // when 2 PAs, equals 2. Otherwise 1

  // - Data Formatter
  wire  [3:0]            crc_loc_stg1;               // one-hot location for the CRC
  wire                   mid_crc_loc_stg1;           // Beat identifier for the mid CRC
  wire                   beat_count_q_is_10;         // Just might be the location of the mid-crc

  wire                   upper_valid_stg1;           // Data valid signal after reordering for AXI
  wire                   lower_valid_stg1;           // Data valid signal after reordering for AXI
  wire                   lower_padded_stg1;          // when 1, the lower word is pad at the end of a packet
  wire                   first_beat_stg1;            // first beat of a packet
  wire [63:0]            ordered_rx_data_stg1;       // Receive data, reordered for AXI
  wire [63:0]            masked_rx_data_stg1;        // Receive data, reordered for AXI, masked AckID for CRC check
  wire                   data_vld_stg1;              // combined data_vld signal - at least one word is valid
  wire                   data_stream_enable_stg1;    // stream enable for both RT and CT
  wire                   control_sym_in_error_cond_cmb; // 11/20/2014
  wire                   not_in_retry_stopped_state; // for CR 825487
  wire                   idle_seq_in_error_cond_cmb;
  wire                   lreq_pd_error;              // this signal detects the PD errors in the LREQ
  wire [1:0]             lreq_reset_dev;             // 12/8/2014
  wire                   in_error_stopped_state;     // Added to fix the CR# 837481, // 12/23/2014
  wire [1:0]             pa_detect_stg0; // 2/5/2015
  // Pipeline stage 2 signals
  // - Carryover from Stage 1
  wire                   framing_end_stg2;           // used with in_packet to indicate the end of a packet
  wire                   framing_start_stg2;         // used with in_packet to indicate the start of a packet
  wire  [3:0]            crc_loc_stg2;               // one-hot location for the CRC
  wire                   dest_dsc_stg2;              // Determination for destination discontinue
  wire                   err_recovery;
  wire                   carryover_stg2;
  wire [1:0]             data_vld_stg0_d;
  wire                   mid_crc_loc_stg2;           // Beat identifier for the mid CRC
  wire                   pr_port_stat_ok;            // Port Status is OK
  wire                   idle2_7_4_beat_err_cmb;     // 2/23/2015, CR # 849824
  // - Input Error Handler - FSM
  wire                   rt_stream_enable_stg2;      // Used to enable the stream for RT

  // - Error Detection Block
  wire                   prx_out_fatal_detect;       // Detected a fatal output error condition
  wire                   prx_force_send_lreq;        // Forces the OLLM TX to send a LREQ
  wire                   prx_out_recoverable_detect; // Detected a recoverable output error
  wire                   prx_in_recoverable_detect;  // Detected a recoverable input error
  wire                   prx_in_retry_detect;        // Detected an input retry event
  wire  [3:0]            prx_cs_crc_check_fail;      // used to generate cs_crc_in_error_cond
  wire                   prx_cs_in_error_cond;       // control symbol error condition detected
  wire                   prx_rcvd_bad_status;        // Detected a bad status control symbol
  wire                   idle2_sync_char_stg0;       // used to indicate sync characters in IDLE2 cases // 11/9/2014
  wire                   in_retry_stopped_state;     // used to indicate Input retry stopped state
  // debug signals
  wire [31:0]            prx_debug;                  // debug signals from the error block
  wire [31:0]            prd_debug;                  // debug signals from the datapath block
  wire                  PR_input_status_good;       // OLLM RX is currently in Output Retry Stopped State
  assign PR_debug = {prx_debug, prd_debug};


  // }}} End wire declarations ------------


  // {{{ Reset Structure ------------------

  // by rule, we must register the resets before we use them. This is not a
  // synchronizing circuit but rather a method to reduce fanout on the resets.
  always @(posedge phy_clk or posedge phy_rst) begin
    if (phy_rst)
      phy_rst_q <= #TCQ 1'b1;
    else
      phy_rst_q <= #TCQ 1'b0;
  end
  always @(posedge log_clk or posedge log_rst) begin
    if (log_rst)
      log_rst_q <= #TCQ 1'b1;
    else
      log_rst_q <= #TCQ 1'b0;
  end

  // }}} End of Reset Structure -----------


  // {{{ OLLM RX CS Decode ------------------
  srio_gen2_v4_1_16_ollm_rx_cs_decode
   #(.TCQ                         (TCQ))
   ollm_rx_cs_decode_inst
    (.phy_clk                     (phy_clk),
    .phy_rst_q                    (phy_rst_q),

    .PP_rx_data                   (PP_rx_data),
    .PP_rx_charisk                (PP_rx_charisk),
    .PP_rx_valid                  (PP_rx_valid),
    .PP_idle2_selected            (PP_idle2_selected),
    .PP_port_initialized          (PP_port_initialized),
    .PR_link_initialized          (PR_link_initialized),

    .PRD_rx_data                  (prd_rx_data),
    .PRD_rx_charisk               (prd_rx_charisk),
    .PRD_rx_valid                 (prd_rx_valid),
    .PRD_idle2_selected           (prd_idle2_selected),
    .PRD_cs_decode                (prd_cs_decode),
    .idle2_sync_char_stg0         (idle2_sync_char_stg0)
    );
  // }}} End of OLLM RX CS Decode ---------


  // {{{ OLLM RX Datapath -------------------
  srio_gen2_v4_1_16_ollm_rx_datapath
   #(.TCQ                         (TCQ),
     .IDLE1                       (IDLE1),
     .IDLE2                       (IDLE2),
     .VC                          (VC),
     .SWITCH_MODE                 (SWITCH_MODE),
     .RETRY                       (RETRY),
     .TARGET_DS                   (TARGET_DS),
     .VC1_CT                      (VC1_CT))
   ollm_rx_datapath_inst
    (.phy_clk                     (phy_clk),
    .phy_rst_q                    (phy_rst_q),
    .PR_phy_rcvd_link_reset       (PR_phy_rcvd_link_reset),
    .prd_debug                    (prd_debug),

    .PRD_rx_data                  (prd_rx_data),
    .PRD_rx_charisk               (prd_rx_charisk),
    .PRD_rx_valid                 (prd_rx_valid),
    .PRD_cs_decode                (prd_cs_decode),
    .PRD_idle2_selected           (prd_idle2_selected),
    .PP_out_of_sync               (PP_out_of_sync),
    .PP_port_initialized          (PP_port_initialized),

    .PR_phyr_tvalid               (PR_phyr_tvalid),
    .BR_phyr_tready               (BR_phyr_tready),
    .PR_phyr_tdata                (PR_phyr_tdata),
    .PR_phyr_tkeep                (PR_phyr_tkeep),
    .PR_phyr_tlast                (PR_phyr_tlast),
    .PR_phyr_tuser                (PR_phyr_tuser),
    .BR_phy_buf_stat              (BR_phy_buf_stat),

    .PT_sent_init_cs              (PT_sent_init_cs),
    .PR_link_initialized          (PR_link_initialized),
    .PR_rewind                    (PR_rewind),
    .PR_phy_rcvd_buf_stat         (PR_phy_rcvd_buf_stat),
    .PR_send_rfr                  (PR_send_rfr),
    .PT_rfr_sent                  (PT_rfr_sent),
    .PR_send_lreq                 (PR_send_lreq),
    .PT_lreq_sent                 (PT_lreq_sent),
    .PR_send_pna                  (PR_send_pna),
    .PT_pna_sent                  (PT_pna_sent),
    .PR_send_pr                   (PR_send_pr),
    .PT_pr_sent                   (PT_pr_sent),
    .PR_send_lresp                (PR_send_lresp),
    .PT_lresp_sent                (PT_lresp_sent),
    .PR_port_stat                 (PR_port_stat),
    .PR_port_stat_ok              (pr_port_stat_ok),
    .PR_output_retry_stop         (PR_output_retry_stop),
    .PR_output_error_stop         (PR_output_error_stop),
    .PR_port_error                (PR_port_error),
    .PR_input_retry_stop          (PR_input_retry_stop),
    .PR_input_error_stop          (PR_input_error_stop),
    .PR_input_status_good         (PR_input_status_good),
    .PR_rcvd_error_free_status    (PR_rcvd_error_free_status),

    .PC_load_ackids               (PC_load_ackids),
    .PC_clr_port_error            (PC_clr_port_error),
    .PC_error_disable             (PC_error_disable),
    .PC_vc_ct                     (PC_vc_ct),
    .PC_vc_en                     (PC_vc_en),
    .PR_rcvd_lresp                (PR_rcvd_lresp),
    .PR_ackid_status              (PR_ackid_status),
    .PR_rcvd_port_stat            (PR_rcvd_port_stat),
    .PR_rcvd_pa_or_pna            (PR_rcvd_pa_or_pna),


    // NOTE - these signals only travel between the sibling modules
    // internal datapath outputs
    // stage 0 inputs (control symbol checking)
    .pd_flag_stg0                (pd_flag_stg0),
    .sc_flag_stg0                (sc_flag_stg0),
    .in_packet_stg0              (in_packet_stg0),
    .sop                         (sop),
    .stomp                       (stomp),
    .eop                         (eop),
    .rfr                         (rfr),
    .lreq                        (lreq),
    .stat                        (stat),
    .mce                         (mce),
    // stage 1 inputs (packet CRC checking)
    .masked_rx_data_stg1         (masked_rx_data_stg1),
    .ordered_rx_data_stg1        (ordered_rx_data_stg1),
    .data_vld_stg1               (data_vld_stg1),
    .data_stream_enable_stg1     (data_stream_enable_stg1),
    .pp_out_of_sync_stg1         (pp_out_of_sync_stg1),
    .pp_port_initialized_stg1    (pp_port_initialized_stg1),
    .crc_loc_stg1                (crc_loc_stg1),
    .mid_crc_loc_stg1            (mid_crc_loc_stg1),
    .beat_count_q_is_10          (beat_count_q_is_10),
    .framing_end_stg1            (framing_end_stg1),
    .framing_start_stg1          (framing_start_stg1),
    .framing_dsc_stg1            (framing_dsc_stg1),
    .upper_valid_stg1            (upper_valid_stg1),
    .lower_valid_stg1            (lower_valid_stg1),
    .lower_padded_stg1           (lower_padded_stg1),
    .first_beat_stg1             (first_beat_stg1),
    .stomp_detect_stg1           (stomp_detect_stg1),
    .lreq_detect_stg1            (lreq_detect_stg1),
    .lreq_in_stat_detect_stg1    (lreq_in_stat_detect_stg1),
    .lresp_detect_stg2           (lresp_detect_stg2),
    .pa_detect_stg1              (pa_detect_stg1),
    .pr_detect_stg1              (pr_detect_stg1),
    .rfr_detect_stg1             (rfr_detect_stg1),
    .pa_ackid_stg1               (pa_ackid_stg1),
    .pr_ackid_stg1               (pr_ackid_stg1),
    .expected_ackid_coef_stg1    (expected_ackid_coef_stg1),
    // stage 2 inputs
    .framing_end_stg2            (framing_end_stg2),
    .framing_start_stg2          (framing_start_stg2),
    .crc_loc_stg2                (crc_loc_stg2),
    .mid_crc_loc_stg2            (mid_crc_loc_stg2),
    .rt_stream_enable_stg2       (rt_stream_enable_stg2),
    .dest_dsc_stg2               (dest_dsc_stg2),
    .err_recovery                (err_recovery),
    .carryover_stg2              (carryover_stg2),
    .data_vld_stg0_d             (data_vld_stg0_d),

    // inputs consumed by datapath
    .prx_out_fatal_detect        (prx_out_fatal_detect),
    .prx_force_send_lreq         (prx_force_send_lreq),
    .prx_out_recoverable_detect  (prx_out_recoverable_detect),
    .prx_in_recoverable_detect   (prx_in_recoverable_detect),
    .prx_in_retry_detect         (prx_in_retry_detect),
    .prx_cs_crc_check_fail       (prx_cs_crc_check_fail),
    .prx_cs_in_error_cond        (prx_cs_in_error_cond),
    .prx_rcvd_bad_status         (prx_rcvd_bad_status),
    .in_retry_stopped_state      (in_retry_stopped_state), // 11/11/2014
    .idle2_sync_char_stg0        (idle2_sync_char_stg0),
    .control_sym_in_error_cond_cmb (control_sym_in_error_cond_cmb),//11/20/2014
    .not_in_retry_stopped_state  (not_in_retry_stopped_state), // 11/25/2014
    .idle_seq_in_error_cond_cmb  (idle_seq_in_error_cond_cmb), // 11/25/2014
    .lreq_pd_error               (lreq_pd_error),
    .lreq_reset_dev              (lreq_reset_dev),// 12/8/2014
    .in_error_stopped_state      (in_error_stopped_state),//12/23/2014
    .pa_detect_stg0              (pa_detect_stg0),// 2/5/2015
    .idle2_7_4_beat_err_cmb      (idle2_7_4_beat_err_cmb) // 2/23/2015, CR # 849824
    );
  // }}} End of OLLM RX Datapath ----------


  // {{{ Error Detection Block --------------
  srio_gen2_v4_1_16_ollm_rx_err_detect
   #(.TCQ                        (TCQ),
     .IDLE1                      (IDLE1),
     .IDLE2                      (IDLE2),
     .MODE_XG                    (MODE_XG),
     .VC                         (VC),
     .SWITCH_MODE                (SWITCH_MODE),
     .RETRY                      (RETRY),
     .LINK_REQUESTS              (LINK_REQUESTS),
     .LINK_WIDTH                (LINK_WIDTH))

   ollm_rx_err_detect_inst
    (.phy_clk                    (phy_clk),
    .phy_rst_q                   (phy_rst_q),
    .log_clk                     (log_clk),
    .log_rst_q                   (log_rst_q),
    .gt_pcs_clk                  (gt_pcs_clk),

    // external inputs
    .PRD_rx_data                 (prd_rx_data),
    .PRD_rx_charisk              (prd_rx_charisk),
    .PRD_idle2_selected          (prd_idle2_selected),
    .PP_gt_decode_error          (PP_gt_decode_error),
    .PP_mode_1x                  (PP_mode_1x), // // updated to fix CR# 835498

    .PR_phyr_tvalid              (PR_phyr_tvalid),
    .BR_phyr_tready              (BR_phyr_tready),
    .PR_phyr_tlast               (PR_phyr_tlast),
    .PR_phyr_tuser               (PR_phyr_tuser),
    .PR_port_stat                (PR_port_stat),
    .PR_port_stat_ok             (pr_port_stat_ok),
    .PR_link_initialized         (PR_link_initialized),
    .PT_sample_next_fm           (PT_sample_next_fm),

    .BR_phy_buf_stat             (BR_phy_buf_stat),
    .PC_next_rcvd_pkt            (PC_next_rcvd_pkt),
    .PC_last_ack                 (PC_last_ack),
    .PC_load_ackids              (PC_load_ackids),
    .PC_load_nextpkt             (PC_load_nextpkt),
    .PC_send_lreq                (PC_send_lreq),
    .PC_lreq_cmd                 (PC_lreq_cmd),
    .PC_link_timeout             (PC_link_timeout),
    .PC_input_maint_only         (PC_input_maint_only),
    .PT_phy_next_fm              (PT_phy_next_fm),
    .PR_output_error_stop        (PR_output_error_stop),
    .PR_output_retry_stop        (PR_output_retry_stop),
    .PR_input_status_good        (PR_input_status_good),
    .PR_send_pna                 (PR_send_pna),
    .PR_send_lreq                (PR_send_lreq),
    .PT_lreq_sent                (PT_lreq_sent),
    .PR_ackid_status             (PR_ackid_status),

    // external outputs
    .PRX_cause                   (PR_cause),
    .PRX_phy_last_ack            (PR_phy_last_ack),
    .PRX_last_good_pkt           (PR_last_good_pkt),
    .PRX_next_rcvd_pkt           (PR_next_rcvd_pkt),
    .PRX_phy_rcvd_mce            (PR_phy_rcvd_mce),
    .prx_debug                   (prx_debug),


    // NOTE - these signals only travel between the sibling modules
    // internal datapath inputs
    // stage 0 inputs (control symbol checking)
    .pd_flag_stg0                (pd_flag_stg0),
    .sc_flag_stg0                (sc_flag_stg0),
    .in_packet_stg0              (in_packet_stg0),
    .sop                         (sop),
    .stomp                       (stomp),
    .eop                         (eop),
    .rfr                         (rfr),
    .lreq                        (lreq),
    .stat                        (stat),
    .mce                         (mce),
    // stage 1 inputs (packet CRC checking)
    .masked_rx_data_stg1         (masked_rx_data_stg1),
    .ordered_rx_data_stg1        (ordered_rx_data_stg1),
    .data_vld_stg1               (data_vld_stg1),
    .data_stream_enable_stg1     (data_stream_enable_stg1),
    .pp_out_of_sync_stg1         (pp_out_of_sync_stg1),
    .pp_port_initialized_stg1    (pp_port_initialized_stg1),
    .crc_loc_stg1                (crc_loc_stg1),
    .mid_crc_loc_stg1            (mid_crc_loc_stg1),
    .beat_count_q_is_10          (beat_count_q_is_10),
    .framing_end_stg1            (framing_end_stg1),
    .framing_start_stg1          (framing_start_stg1),
    .framing_dsc_stg1            (framing_dsc_stg1),
    .upper_valid_stg1            (upper_valid_stg1),
    .lower_valid_stg1            (lower_valid_stg1),
    .lower_padded_stg1           (lower_padded_stg1),
    .first_beat_stg1             (first_beat_stg1),
    .stomp_detect_stg1           (stomp_detect_stg1),
    .lreq_detect_stg1            (lreq_detect_stg1),
    .lreq_in_stat_detect_stg1    (lreq_in_stat_detect_stg1),
    .lresp_detect_stg2           (lresp_detect_stg2),
    .pa_detect_stg1              (pa_detect_stg1),
    .pr_detect_stg1              (pr_detect_stg1),
    .rfr_detect_stg1             (rfr_detect_stg1),
    .pa_ackid_stg1               (pa_ackid_stg1),
    .pr_ackid_stg1               (pr_ackid_stg1),
    .expected_ackid_coef_stg1    (expected_ackid_coef_stg1),
    // stage 2 inputs
    .framing_end_stg2            (framing_end_stg2),
    .framing_start_stg2          (framing_start_stg2),
    .crc_loc_stg2                (crc_loc_stg2),
    .mid_crc_loc_stg2            (mid_crc_loc_stg2),
    .rt_stream_enable_stg2       (rt_stream_enable_stg2),
    .dest_dsc_stg2               (dest_dsc_stg2),
    .err_recovery                (err_recovery),
    .carryover_stg2              (carryover_stg2),
    .data_vld_stg0_d             (data_vld_stg0_d),

    // outputs consumed by datapath
    .prx_out_fatal_detect        (prx_out_fatal_detect),
    .prx_force_send_lreq         (prx_force_send_lreq),
    .prx_out_recoverable_detect  (prx_out_recoverable_detect),
    .prx_in_recoverable_detect   (prx_in_recoverable_detect),
    .prx_in_retry_detect         (prx_in_retry_detect),
    .prx_cs_crc_check_fail       (prx_cs_crc_check_fail),
    .prx_cs_in_error_cond        (prx_cs_in_error_cond),
    .prx_rcvd_bad_status         (prx_rcvd_bad_status),
    .idle2_sync_char_stg0        (idle2_sync_char_stg0),           //11/9/2014
    .in_retry_stopped_state      (in_retry_stopped_state),         // 11/11/2014
    .control_sym_in_error_cond_cmb (control_sym_in_error_cond_cmb), //11/20/2014
    .not_in_retry_stopped_state  (not_in_retry_stopped_state), // 11/25/2014
    .idle_seq_in_error_cond_cmb  (idle_seq_in_error_cond_cmb), // 11/25/2014
    .lreq_pd_error               (lreq_pd_error),
    .lreq_reset_dev              (lreq_reset_dev),// 12/8/2014
    .in_error_stopped_state      (in_error_stopped_state),//12/23/2014
    .pa_detect_stg0              (pa_detect_stg0), //2/5/2015
    .idle2_7_4_beat_err_cmb      (idle2_7_4_beat_err_cmb) // 2/23/2015, CR # 849824
    );
  // }}} End of Error Detection Block -----

endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
//
// CRC5_20
//
// Description:
// This module calculates the 5-bit CRC for 20-bits in a short control 
// symbol.This was taken from section 3.6.2 CRC generation, Table 3-9 in 
// the PHY layer Spec.
//
// REQ: req_pt_short_cs_polynomial
// REQ: req_pt_crc5_init_value
// ---------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_crc5_20
  (
    input       [0:18]  din,   // Data 
    output wire [0:4]   crc    // Calculated CRC-5     
  );

  assign crc[0] = din[18]  ^ din[16] ^ din[15] ^ din[12] ^ din[10] ^ din[5]  ^ 
                  din[4]   ^ din[3]  ^ din[1]  ^ din[0];

  assign crc[1] = !din[18] ^ din[17] ^ din[15] ^ din[13] ^ din[12] ^ din[11] ^
                   din[10] ^ din[6]  ^ din[3]  ^ din[2]  ^ din[0];

  assign crc[2] = !din[18] ^ din[16] ^ din[14] ^ din[13] ^ din[12] ^ din[11] ^
                   din[7]  ^ din[4]  ^ din[3]  ^ din[1];

  assign crc[3] = !din[18] ^ din[17] ^ din[16] ^ din[14] ^ din[13] ^ din[10] ^
                   din[8]  ^ din[3]  ^ din[2]  ^ din[1];

  assign crc[4] = din[18]  ^ din[17] ^ din[15] ^ din[14] ^ din[11] ^ din[9]  ^
                  din[4]   ^ din[3]  ^ din[2]  ^ din[0];

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//-------------------------------------------------------------------------
// CRC16_16
//
// Description:
// This module takes 48-bits of data and a 16-bit CRC to produce a new CRC
//
// REQ: req_pt_crc16_polynomial
//
// IPCV - easics used
// Equations obtained from: 
// http://www.easics.be/webtools/crctool
// ------------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_crc16_48
  ( 
    input       [47:0] din,   // Input Data
    input       [15:0] cin,   // Input CRC
    output wire [15:0] crc    // New Output CRC
  );

  assign crc[0]  = din[42] ^ din[35] ^ din[33] ^ din[32] ^ din[28] ^ din[27] ^ din[26] ^ 
                   din[22] ^ din[20] ^ din[19] ^ din[12] ^ din[11] ^ din[8]  ^ din[4]  ^ 
                   din[0]  ^ cin[0]  ^ cin[1]  ^ cin[3]  ^ cin[10];

  assign crc[1]  = din[43] ^ din[36] ^ din[34] ^ din[33] ^ din[29] ^ din[28] ^ din[27] ^ 
                   din[23] ^ din[21] ^ din[20] ^ din[13] ^ din[12] ^ din[9]  ^ din[5]  ^ 
                   din[1]  ^ cin[1]  ^ cin[2]  ^ cin[4]  ^ cin[11];

  assign crc[2]  = din[44] ^ din[37] ^ din[35] ^ din[34] ^ din[30] ^ din[29] ^ din[28] ^ 
                   din[24] ^ din[22] ^ din[21] ^ din[14] ^ din[13] ^ din[10] ^ din[6]  ^ 
                   din[2]  ^ cin[2]  ^ cin[3]  ^ cin[5]  ^ cin[12];

  assign crc[3]  = din[45] ^ din[38] ^ din[36] ^ din[35] ^ din[31] ^ din[30] ^ din[29] ^ 
                   din[25] ^ din[23] ^ din[22] ^ din[15] ^ din[14] ^ din[11] ^ din[7]  ^ 
                   din[3]  ^ cin[3]  ^ cin[4]  ^ cin[6]  ^ cin[13];

  assign crc[4]  = din[46] ^ din[39] ^ din[37] ^ din[36] ^ din[32] ^ din[31] ^ din[30] ^ 
                   din[26] ^ din[24] ^ din[23] ^ din[16] ^ din[15] ^ din[12] ^ din[8]  ^ 
                   din[4]  ^ cin[0]  ^ cin[4]  ^ cin[5]  ^ cin[7]  ^ cin[14];

  assign crc[5]  = din[47] ^ din[42] ^ din[40] ^ din[38] ^ din[37] ^ din[35] ^ din[31] ^ 
                   din[28] ^ din[26] ^ din[25] ^ din[24] ^ din[22] ^ din[20] ^ din[19] ^ 
                   din[17] ^ din[16] ^ din[13] ^ din[12] ^ din[11] ^ din[9]  ^ din[8]  ^ 
                   din[5]  ^ din[4]  ^ din[0]  ^ cin[3]  ^ cin[5]  ^ cin[6]  ^ cin[8]  ^ 
                   cin[10] ^ cin[15];

  assign crc[6]  = din[43] ^ din[41] ^ din[39] ^ din[38] ^ din[36] ^ din[32] ^ din[29] ^ 
                   din[27] ^ din[26] ^ din[25] ^ din[23] ^ din[21] ^ din[20] ^ din[18] ^ 
                   din[17] ^ din[14] ^ din[13] ^ din[12] ^ din[10] ^ din[9]  ^ din[6] ^ 
                   din[5]  ^ din[1]  ^ cin[0]  ^ cin[4]  ^ cin[6]  ^ cin[7]  ^ cin[9] ^ 
                   cin[11];

  assign crc[7]  = din[44] ^ din[42] ^ din[40] ^ din[39] ^ din[37] ^ din[33] ^ din[30] ^ 
                   din[28] ^ din[27] ^ din[26] ^ din[24] ^ din[22] ^ din[21] ^ din[19] ^ 
                   din[18] ^ din[15] ^ din[14] ^ din[13] ^ din[11] ^ din[10] ^ din[7]  ^ 
                   din[6]  ^ din[2]  ^ cin[1]  ^ cin[5]  ^ cin[7]  ^ cin[8]  ^ cin[10] ^ 
                   cin[12];

  assign crc[8]  = din[45] ^ din[43] ^ din[41] ^ din[40] ^ din[38] ^ din[34] ^ din[31] ^ 
                   din[29] ^ din[28] ^ din[27] ^ din[25] ^ din[23] ^ din[22] ^ din[20] ^ 
                   din[19] ^ din[16] ^ din[15] ^ din[14] ^ din[12] ^ din[11] ^ din[8]  ^ 
                   din[7]  ^ din[3]  ^ cin[2]  ^ cin[6]  ^ cin[8]  ^ cin[9]  ^ cin[11] ^ 
                   cin[13];
  assign crc[9]  = din[46] ^ din[44] ^ din[42] ^ din[41] ^ din[39] ^ din[35] ^ din[32] ^ 
                   din[30] ^ din[29] ^ din[28] ^ din[26] ^ din[24] ^ din[23] ^ din[21] ^ 
                   din[20] ^ din[17] ^ din[16] ^ din[15] ^ din[13] ^ din[12] ^ din[9]  ^ 
                   din[8]  ^ din[4]  ^ cin[0]  ^ cin[3]  ^ cin[7]  ^ cin[9]  ^ cin[10] ^ 
                   cin[12] ^ cin[14];
  assign crc[10] = din[47] ^ din[45] ^ din[43] ^ din[42] ^ din[40] ^ din[36] ^ din[33] ^ 
                   din[31] ^ din[30] ^ din[29] ^ din[27] ^ din[25] ^ din[24] ^ din[22] ^ 
                   din[21] ^ din[18] ^ din[17] ^ din[16] ^ din[14] ^ din[13] ^ din[10] ^ 
                   din[9]  ^ din[5]  ^ cin[1]  ^ cin[4]  ^ cin[8]  ^ cin[10] ^ cin[11] ^ 
                   cin[13] ^ cin[15];
  assign crc[11] = din[46] ^ din[44] ^ din[43] ^ din[41] ^ din[37] ^ din[34] ^ din[32] ^ 
                   din[31] ^ din[30] ^ din[28] ^ din[26] ^ din[25] ^ din[23] ^ din[22] ^ 
                   din[19] ^ din[18] ^ din[17] ^ din[15] ^ din[14] ^ din[11] ^ din[10] ^ 
                   din[6]  ^ cin[0]  ^ cin[2]  ^ cin[5]  ^ cin[9]  ^ cin[11] ^ cin[12] ^ 
                   cin[14];
  assign crc[12] = din[47] ^ din[45] ^ din[44] ^ din[38] ^ din[31] ^ din[29] ^ din[28] ^ 
                   din[24] ^ din[23] ^ din[22] ^ din[18] ^ din[16] ^ din[15] ^ din[8]  ^ 
                   din[7]  ^ din[4]  ^ din[0]  ^ cin[6]  ^ cin[12] ^ cin[13] ^ cin[15];
  assign crc[13] = din[46] ^ din[45] ^ din[39] ^ din[32] ^ din[30] ^ din[29] ^ din[25] ^ 
                   din[24] ^ din[23] ^ din[19] ^ din[17] ^ din[16] ^ din[9]  ^ din[8]  ^ 
                   din[5]  ^ din[1]  ^ cin[0]  ^ cin[7]  ^ cin[13] ^ cin[14];
  assign crc[14] = din[47] ^ din[46] ^ din[40] ^ din[33] ^ din[31] ^ din[30] ^ din[26] ^ 
                   din[25] ^ din[24] ^ din[20] ^ din[18] ^ din[17] ^ din[10] ^ din[9]  ^ 
                   din[6]  ^ din[2]  ^ cin[1]  ^ cin[8]  ^ cin[14] ^ cin[15];
  assign crc[15] = din[47] ^ din[41] ^ din[34] ^ din[32] ^ din[31] ^ din[27] ^ din[26] ^ 
                   din[25] ^ din[21] ^ din[19] ^ din[18] ^ din[11] ^ din[10] ^ din[7]  ^ 
                   din[3]  ^ cin[0]  ^ cin[2]  ^ cin[9]  ^ cin[15];

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
//
// CRC13_35
//
// Description:
// This module calculates the 13-bit CRC for the 34-bits in a long control 
// symbol. These equations were derived from section 3.6.4 CRC-13 Parallel Code
// Generation, Table 3-10 of the PHY layer spec.
// 
// REQ: req_pt_long_cs_polynomial
// REQ: req_pt_crc13_init_value
// ---------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_crc13_35
  (
    output wire [0:12]  crc,   // Calculated CRC-13
    input       [0:34]  din    // Data 
  );
 
  assign crc[0]  = din[32] ^ din[30] ^ din[29] ^ din[27] ^ din[26] ^ din[25] ^ din[23] ^
                   din[21] ^ din[19] ^ din[14] ^ din[9]  ^ din[6]  ^ din[4];

  assign crc[1]  = din[33] ^ din[31] ^ din[30] ^ din[28] ^ din[27] ^ din[26] ^ din[24] ^
                   din[22] ^ din[20] ^ din[15] ^ din[10] ^ din[7]  ^ din[5]  ^ din[0];

  assign crc[2]  = din[34] ^ din[32] ^ din[31] ^ din[29] ^ din[28] ^ din[27] ^ din[25] ^
                   din[23] ^ din[21] ^ din[16] ^ din[11] ^ din[8]  ^ din[6]  ^ din[1];

  assign crc[3]  = din[33] ^ din[28] ^ din[27] ^ din[25] ^ din[24] ^ din[23] ^ din[22] ^
                   din[21] ^ din[19] ^ din[17] ^ din[14] ^ din[12] ^ din[7]  ^ din[6]  ^
                   din[4]  ^ din[2];

  assign crc[4]  = din[34] ^ din[29] ^ din[28] ^ din[26] ^ din[25] ^ din[24] ^ din[23] ^
                   din[22] ^ din[20] ^ din[18] ^ din[15] ^ din[13] ^ din[8] ^ din[7]   ^
                   din[5]  ^ din[3];

  assign crc[5]  = din[32] ^ din[24] ^ din[16] ^ din[8] ^ din[0];

  assign crc[6]  = din[33] ^ din[25] ^ din[17] ^ din[9] ^ din[1];

  assign crc[7]  = din[34] ^ din[26] ^ din[18] ^ din[10] ^ din[2];

  assign crc[8]  = din[32] ^ din[30] ^ din[29] ^ din[26] ^ din[25] ^ din[23] ^ din[21] ^
                   din[14] ^ din[11] ^ din[9]  ^ din[6]  ^ din[4]  ^ din[3];

  assign crc[9]  = din[33] ^ din[31] ^ din[30] ^ din[27] ^ din[26] ^ din[24] ^ din[22] ^
                   din[15] ^ din[12] ^ din[10] ^ din[7]  ^ din[5]  ^ din[4]  ^ din[0];

  assign crc[10] = din[34] ^ din[32] ^ din[31] ^ din[28] ^ din[27] ^ din[25] ^ din[23] ^
                   din[16] ^ din[13] ^ din[11] ^ din[8]  ^ din[6]  ^ din[5]  ^ din[1];

  assign crc[11] = din[33] ^ din[30] ^ din[28] ^ din[27] ^ din[25] ^ din[24] ^ din[23] ^
                   din[21] ^ din[19] ^ din[17] ^ din[12] ^ din[7]  ^ din[4]  ^ din[2];

  assign crc[12] = din[34] ^ din[31] ^ din[29] ^ din[28] ^ din[26] ^ din[25] ^ din[24] ^
                   din[22] ^ din[20] ^ din[18] ^ din[13] ^ din[8]  ^ din[5]  ^ din[3];

endmodule
  
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//-------------------------------------------------------------------------
// CRC16_16
//
// Description:
// This module takes 16-bits of data and a 16-bit CRC to produce a new CRC
//
// REQ: req_pt_crc16_polynomial
//
// IPCV - easics used
// Equations obtained from: 
// http://www.easics.be/webtools/crctool
// ------------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_crc16_16
  ( 
    input       [15:0] din,  // Input Data
    input       [15:0] cin,  // Input CRC
    output wire [15:0] crc   // Output new CRC
  );

  assign crc[0]  = din[12] ^ din[11] ^ din[8]  ^ din[4]  ^ din[0]  ^ cin[0]  ^ cin[4]  ^ 
                   cin[8]  ^ cin[11] ^ cin[12];

  assign crc[1]  = din[13] ^ din[12] ^ din[9]  ^ din[5]  ^ din[1]  ^ cin[1]  ^ cin[5]  ^ 
                   cin[9]  ^ cin[12] ^ cin[13];

  assign crc[2]  = din[14] ^ din[13] ^ din[10] ^ din[6]  ^ din[2]  ^ cin[2]  ^ cin[6]  ^ 
                   cin[10] ^ cin[13] ^ cin[14];

  assign crc[3]  = din[15] ^ din[14] ^ din[11] ^ din[7]  ^ din[3]  ^ cin[3]  ^ cin[7]  ^ 
                   cin[11] ^ cin[14] ^ cin[15];

  assign crc[4]  = din[15] ^ din[12] ^ din[8]  ^ din[4]  ^ cin[4]  ^ cin[8]  ^ cin[12] ^ 
                   cin[15];
  assign crc[5]  = din[13] ^ din[12] ^ din[11] ^ din[9]  ^ din[8]  ^ din[5]  ^ din[4]  ^ 
                   din[0]  ^ cin[0]  ^ cin[4]  ^ cin[5]  ^ cin[8]  ^ cin[9]  ^ cin[11] ^ 
                   cin[12] ^ cin[13];

  assign crc[6]  = din[14] ^ din[13] ^ din[12] ^ din[10] ^ din[9]  ^ din[6]  ^ din[5]  ^ 
                   din[1]  ^ cin[1]  ^ cin[5]  ^ cin[6]  ^ cin[9]  ^ cin[10] ^ cin[12] ^ 
                   cin[13] ^ cin[14];

  assign crc[7]  = din[15] ^ din[14] ^ din[13] ^ din[11] ^ din[10] ^ din[7]  ^ din[6]  ^ 
                   din[2]  ^ cin[2]  ^ cin[6]  ^ cin[7]  ^ cin[10] ^ cin[11] ^ cin[13] ^ 
                   cin[14] ^ cin[15];

  assign crc[8]  = din[15] ^ din[14] ^ din[12] ^ din[11] ^ din[8]  ^ din[7]  ^ din[3]  ^ 
                   cin[3]  ^ cin[7]  ^ cin[8]  ^ cin[11] ^ cin[12] ^ cin[14] ^ cin[15];

  assign crc[9]  = din[15] ^ din[13] ^ din[12] ^ din[9]  ^ din[8]  ^ din[4]  ^ cin[4]  ^ 
                   cin[8]  ^ cin[9]  ^ cin[12] ^ cin[13] ^ cin[15];

  assign crc[10] = din[14] ^ din[13] ^ din[10] ^ din[9]  ^ din[5]  ^ cin[5]  ^ cin[9]  ^ 
                   cin[10] ^ cin[13] ^ cin[14];

  assign crc[11] = din[15] ^ din[14] ^ din[11] ^ din[10] ^ din[6]  ^ cin[6]  ^ cin[10] ^ 
                   cin[11] ^ cin[14] ^ cin[15];

  assign crc[12] = din[15] ^ din[8]  ^ din[7]  ^ din[4]  ^ din[0]  ^ cin[0]  ^ cin[4]  ^ 
                   cin[7] ^ cin[8]  ^ cin[15];

  assign crc[13] = din[9]  ^ din[8]  ^ din[5]  ^ din[1]  ^ cin[1]  ^ cin[5]  ^ cin[8]  ^ 
                   cin[9];

  assign crc[14] = din[10] ^ din[9]  ^ din[6]  ^ din[2]  ^ cin[2]  ^ cin[6]  ^ cin[9]  ^
                   cin[10];

  assign crc[15] = din[11] ^ din[10] ^ din[7]  ^ din[3]  ^ cin[3]  ^ cin[7]  ^ cin[10] ^ 
                   cin[11];

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//-------------------------------------------------------------------------
// CRC16_64
//
// Description:
// This module takes 64-bits of data and a 16-bit CRC to produce a new CRC
//
// REQ: req_pt_crc16_polynomial
//
// IPCV - easics used
// Equations obtained from: 
// http://www.easics.be/webtools/crctool
// ------------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_crc16_64
  ( 
    input  [63:0] din,  // Input Data
    input  [15:0] cin,  // Input CRC
    output [15:0] crc   // New output CRC
  );

  assign crc[0]  = din[63] ^ din[58] ^ din[56] ^ din[55] ^ din[52] ^ din[51] ^ din[49] ^ 
                   din[48] ^ din[42] ^ din[35] ^ din[33] ^ din[32] ^ din[28] ^ din[27] ^ 
                   din[26] ^ din[22] ^ din[20] ^ din[19] ^ din[12] ^ din[11] ^ din[8]  ^ 
                   din[4]  ^ din[0]  ^ cin[0]  ^ cin[1]  ^ cin[3]  ^ cin[4]  ^ cin[7]  ^ 
                   cin[8]  ^ cin[10] ^ cin[15];

  assign crc[1]  = din[59] ^ din[57] ^ din[56] ^ din[53] ^ din[52] ^ din[50] ^ din[49] ^ 
                   din[43] ^ din[36] ^ din[34] ^ din[33] ^ din[29] ^ din[28] ^ din[27] ^ 
                   din[23] ^ din[21] ^ din[20] ^ din[13] ^ din[12] ^ din[9]  ^ din[5]  ^ 
                   din[1]  ^ cin[1]  ^ cin[2]  ^ cin[4]  ^ cin[5]  ^ cin[8]  ^ cin[9]  ^ 
                   cin[11];

  assign crc[2]  = din[60] ^ din[58] ^ din[57] ^ din[54] ^ din[53] ^ din[51] ^ din[50] ^ 
                   din[44] ^ din[37] ^ din[35] ^ din[34] ^ din[30] ^ din[29] ^ din[28] ^ 
                   din[24] ^ din[22] ^ din[21] ^ din[14] ^ din[13] ^ din[10] ^ din[6]  ^ 
                   din[2]  ^ cin[2]  ^ cin[3]  ^ cin[5]  ^ cin[6]  ^ cin[9]  ^ cin[10] ^ 
                   cin[12];
  assign crc[3]  = din[61] ^ din[59] ^ din[58] ^ din[55] ^ din[54] ^ din[52] ^ din[51] ^ 
                   din[45] ^ din[38] ^ din[36] ^ din[35] ^ din[31] ^ din[30] ^ din[29] ^ 
                   din[25] ^ din[23] ^ din[22] ^ din[15] ^ din[14] ^ din[11] ^ din[7]  ^ 
                   din[3]  ^ cin[3]  ^ cin[4]  ^ cin[6]  ^ cin[7]  ^ cin[10] ^ cin[11] ^ 
                   cin[13];

  assign crc[4]  = din[62] ^ din[60] ^ din[59] ^ din[56] ^ din[55] ^ din[53] ^ din[52] ^ 
                   din[46] ^ din[39] ^ din[37] ^ din[36] ^ din[32] ^ din[31] ^ din[30] ^ 
                   din[26] ^ din[24] ^ din[23] ^ din[16] ^ din[15] ^ din[12] ^ din[8]  ^ 
                   din[4]  ^ cin[4]  ^ cin[5]  ^ cin[7]  ^ cin[8]  ^ cin[11] ^ cin[12] ^ 
                   cin[14];

  assign crc[5]  = din[61] ^ din[60] ^ din[58] ^ din[57] ^ din[55] ^ din[54] ^ din[53] ^ 
                   din[52] ^ din[51] ^ din[49] ^ din[48] ^ din[47] ^ din[42] ^ din[40] ^ 
                   din[38] ^ din[37] ^ din[35] ^ din[31] ^ din[28] ^ din[26] ^ din[25] ^ 
                   din[24] ^ din[22] ^ din[20] ^ din[19] ^ din[17] ^ din[16] ^ din[13] ^ 
                   din[12] ^ din[11] ^ din[9]  ^ din[8]  ^ din[5]  ^ din[4]  ^ din[0]  ^ 
                   cin[0]  ^ cin[1]  ^ cin[3]  ^ cin[4]  ^ cin[5]  ^ cin[6]  ^ cin[7]  ^ 
                   cin[9]  ^ cin[10] ^ cin[12] ^ cin[13];

  assign crc[6]  = din[62] ^ din[61] ^ din[59] ^ din[58] ^ din[56] ^ din[55] ^ din[54] ^ 
                   din[53] ^ din[52] ^ din[50] ^ din[49] ^ din[48] ^ din[43] ^ din[41] ^ 
                   din[39] ^ din[38] ^ din[36] ^ din[32] ^ din[29] ^ din[27] ^ din[26] ^ 
                   din[25] ^ din[23] ^ din[21] ^ din[20] ^ din[18] ^ din[17] ^ din[14] ^ 
                   din[13] ^ din[12] ^ din[10] ^ din[9]  ^ din[6]  ^ din[5]  ^ din[1]  ^ 
                   cin[0]  ^ cin[1]  ^ cin[2]  ^ cin[4]  ^ cin[5]  ^ cin[6]  ^ cin[7]  ^ 
                   cin[8]  ^ cin[10] ^ cin[11] ^ cin[13] ^ cin[14];

  assign crc[7]  = din[63] ^ din[62] ^ din[60] ^ din[59] ^ din[57] ^ din[56] ^ din[55] ^ 
                   din[54] ^ din[53] ^ din[51] ^ din[50] ^ din[49] ^ din[44] ^ din[42] ^ 
                   din[40] ^ din[39] ^ din[37] ^ din[33] ^ din[30] ^ din[28] ^ din[27] ^ 
                   din[26] ^ din[24] ^ din[22] ^ din[21] ^ din[19] ^ din[18] ^ din[15] ^ 
                   din[14] ^ din[13] ^ din[11] ^ din[10] ^ din[7]  ^ din[6]  ^ din[2]  ^ 
                   cin[1]  ^ cin[2]  ^ cin[3]  ^ cin[5]  ^ cin[6]  ^ cin[7]  ^ cin[8]  ^ 
                   cin[9]  ^ cin[11] ^ cin[12] ^ cin[14] ^ cin[15];

  assign crc[8]  = din[63] ^ din[61] ^ din[60] ^ din[58] ^ din[57] ^ din[56] ^ din[55] ^ 
                   din[54] ^ din[52] ^ din[51] ^ din[50] ^ din[45] ^ din[43] ^ din[41] ^ 
                   din[40] ^ din[38] ^ din[34] ^ din[31] ^ din[29] ^ din[28] ^ din[27] ^ 
                   din[25] ^ din[23] ^ din[22] ^ din[20] ^ din[19] ^ din[16] ^ din[15] ^ 
                   din[14] ^ din[12] ^ din[11] ^ din[8]  ^ din[7]  ^ din[3]  ^ cin[2]  ^ 
                   cin[3]  ^ cin[4]  ^ cin[6]  ^ cin[7]  ^ cin[8]  ^ cin[9]  ^ cin[10] ^ 
                   cin[12] ^ cin[13] ^ cin[15];

  assign crc[9]  = din[62] ^ din[61] ^ din[59] ^ din[58] ^ din[57] ^ din[56] ^ din[55] ^ 
                   din[53] ^ din[52] ^ din[51] ^ din[46] ^ din[44] ^ din[42] ^ din[41] ^ 
                   din[39] ^ din[35] ^ din[32] ^ din[30] ^ din[29] ^ din[28] ^ din[26] ^ 
                   din[24] ^ din[23] ^ din[21] ^ din[20] ^ din[17] ^ din[16] ^ din[15] ^ 
                   din[13] ^ din[12] ^ din[9]  ^ din[8]  ^ din[4]  ^ cin[3]  ^ cin[4]  ^ 
                   cin[5]  ^ cin[7]  ^ cin[8]  ^ cin[9]  ^ cin[10] ^ cin[11] ^ cin[13] ^ 
                   cin[14];

  assign crc[10] = din[63] ^ din[62] ^ din[60] ^ din[59] ^ din[58] ^ din[57] ^ din[56] ^ 
                   din[54] ^ din[53] ^ din[52] ^ din[47] ^ din[45] ^ din[43] ^ din[42] ^ 
                   din[40] ^ din[36] ^ din[33] ^ din[31] ^ din[30] ^ din[29] ^ din[27] ^ 
                   din[25] ^ din[24] ^ din[22] ^ din[21] ^ din[18] ^ din[17] ^ din[16] ^ 
                   din[14] ^ din[13] ^ din[10] ^ din[9]  ^ din[5]  ^ cin[4]  ^ cin[5]  ^ 
                   cin[6]   ^ cin[8] ^ cin[9]  ^ cin[10] ^ cin[11] ^ cin[12] ^ cin[14] ^ 
                   cin[15];

  assign crc[11] = din[63] ^ din[61] ^ din[60] ^ din[59] ^ din[58] ^ din[57] ^ din[55] ^ 
                   din[54] ^ din[53] ^ din[48] ^ din[46] ^ din[44] ^ din[43] ^ din[41] ^ 
                   din[37] ^ din[34] ^ din[32] ^ din[31] ^ din[30] ^ din[28] ^ din[26] ^ 
                   din[25] ^ din[23] ^ din[22] ^ din[19] ^ din[18] ^ din[17] ^ din[15] ^ 
                   din[14] ^ din[11] ^ din[10] ^ din[6]  ^ cin[0]  ^ cin[5]  ^ cin[6]  ^ 
                   cin[7]  ^ cin[9]  ^ cin[10] ^ cin[11] ^ cin[12] ^ cin[13] ^ cin[15];

  assign crc[12] = din[63] ^ din[62] ^ din[61] ^ din[60] ^ din[59] ^ din[54] ^ din[52] ^ 
                   din[51] ^ din[48] ^ din[47] ^ din[45] ^ din[44] ^ din[38] ^ din[31] ^ 
                   din[29] ^ din[28] ^ din[24] ^ din[23] ^ din[22] ^ din[18] ^ din[16] ^ 
                   din[15] ^ din[8]  ^ din[7]  ^ din[4]  ^ din[0]  ^ cin[0]  ^ cin[3]  ^ 
                   cin[4]  ^ cin[6]  ^ cin[11] ^ cin[12] ^ cin[13] ^ cin[14] ^ cin[15];

  assign crc[13] = din[63] ^ din[62] ^ din[61] ^ din[60] ^ din[55] ^ din[53] ^ din[52] ^ 
                   din[49] ^ din[48] ^ din[46] ^ din[45] ^ din[39] ^ din[32] ^ din[30] ^ 
                   din[29] ^ din[25] ^ din[24] ^ din[23] ^ din[19] ^ din[17] ^ din[16] ^ 
                   din[9]  ^ din[8]  ^ din[5]  ^ din[1]  ^ cin[0]  ^ cin[1]  ^ cin[4]  ^ 
                   cin[5]  ^ cin[7]  ^ cin[12] ^ cin[13] ^ cin[14] ^ cin[15];

  assign crc[14] = din[63] ^ din[62] ^ din[61] ^ din[56] ^ din[54] ^ din[53] ^ din[50] ^ 
                   din[49] ^ din[47] ^ din[46] ^ din[40] ^ din[33] ^ din[31] ^ din[30] ^ 
                   din[26] ^ din[25] ^ din[24] ^ din[20] ^ din[18] ^ din[17] ^ din[10] ^ 
                   din[9]  ^ din[6]  ^ din[2]  ^ cin[1]  ^ cin[2]  ^ cin[5]  ^ cin[6]  ^ 
                   cin[8]  ^ cin[13] ^ cin[14] ^ cin[15];

  assign crc[15] = din[63] ^ din[62] ^ din[57] ^ din[55] ^ din[54] ^ din[51] ^ din[50] ^ 
                   din[48] ^ din[47] ^ din[41] ^ din[34] ^ din[32] ^ din[31] ^ din[27] ^ 
                   din[26] ^ din[25] ^ din[21] ^ din[19] ^ din[18] ^ din[11] ^ din[10] ^ 
                   din[7]  ^ din[3]  ^ cin[0]  ^ cin[2]  ^ cin[3]  ^ cin[6]  ^ cin[7]  ^ 
                   cin[9]  ^ cin[14] ^ cin[15];

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//-------------------------------------------------------------------------
// CRC16_16
//
// Description:
// This module takes 32-bits of data and a 16-bit CRC to produce a new CRC
//
// REQ: req_pt_crc16_polynomial
//
// IPCV - easics used
// Equations obtained from: 
// http://www.easics.be/webtools/crctool
// ------------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_crc16_32
  ( 
    input       [31:0] din, // Input Data
    input       [15:0] cin, // Input CRC
    output wire [15:0] crc  // New Output CRC
  );
 
  assign crc[0]  = din[28] ^ din[27] ^ din[26] ^ din[22] ^ din[20] ^ din[19] ^ din[12] ^ 
                   din[11] ^ din[8]  ^ din[4]  ^ din[0]  ^ cin[3]  ^ cin[4]  ^ cin[6]  ^ 
                   cin[10] ^ cin[11] ^ cin[12];

  assign crc[1]  = din[29] ^ din[28] ^ din[27] ^ din[23] ^ din[21] ^ din[20] ^ din[13] ^ 
                   din[12] ^ din[9]  ^ din[5]  ^ din[1]  ^ cin[4]  ^ cin[5]  ^ cin[7]  ^ 
                   cin[11] ^ cin[12] ^ cin[13];

  assign crc[2]  = din[30] ^ din[29] ^ din[28] ^ din[24] ^ din[22] ^ din[21] ^ din[14] ^ 
                   din[13] ^ din[10] ^ din[6]  ^ din[2]  ^ cin[5]  ^ cin[6]  ^ cin[8]  ^ 
                   cin[12] ^ cin[13] ^ cin[14];

  assign crc[3]  = din[31] ^ din[30] ^ din[29] ^ din[25] ^ din[23] ^ din[22] ^ din[15] ^ 
                   din[14] ^ din[11] ^ din[7]  ^ din[3]  ^ cin[6]  ^ cin[7]  ^ cin[9]  ^ 
                   cin[13] ^ cin[14] ^ cin[15];

  assign crc[4]  = din[31] ^ din[30] ^ din[26] ^ din[24] ^ din[23] ^ din[16] ^ din[15] ^ 
                   din[12] ^ din[8]  ^ din[4]  ^ cin[0]  ^ cin[7]  ^ cin[8]  ^ cin[10] ^ 
                   cin[14] ^ cin[15];

  assign crc[5]  = din[31] ^ din[28] ^ din[26] ^ din[25] ^ din[24] ^ din[22] ^ din[20] ^ 
                   din[19] ^ din[17] ^ din[16] ^ din[13] ^ din[12] ^ din[11] ^ din[9]  ^ 
                   din[8]  ^ din[5]  ^ din[4]  ^ din[0]  ^ cin[0]  ^ cin[1]  ^ cin[3]  ^ 
                   cin[4] ^  cin[6]  ^ cin[8]  ^ cin[9]  ^ cin[10] ^ cin[12] ^ cin[15];

  assign crc[6]  = din[29] ^ din[27] ^ din[26] ^ din[25] ^ din[23] ^ din[21] ^ din[20] ^ 
                   din[18] ^ din[17] ^ din[14] ^ din[13] ^ din[12] ^ din[10] ^ din[9]  ^ 
                   din[6]  ^ din[5]  ^ din[1]  ^ cin[1]  ^ cin[2]  ^ cin[4]  ^ cin[5]  ^ 
                   cin[7] ^  cin[9]  ^ cin[10] ^ cin[11] ^ cin[13];

  assign crc[7]  = din[30] ^ din[28] ^ din[27] ^ din[26] ^ din[24] ^ din[22] ^ din[21] ^ 
                   din[19] ^ din[18] ^ din[15] ^ din[14] ^ din[13] ^ din[11] ^ din[10] ^ 
                   din[7]  ^ din[6]  ^ din[2]  ^ cin[2]  ^ cin[3]  ^ cin[5]  ^ cin[6]  ^ 
                   cin[8]  ^ cin[10] ^ cin[11] ^ cin[12] ^ cin[14];

  assign crc[8]  = din[31] ^ din[29] ^ din[28] ^ din[27] ^ din[25] ^ din[23] ^ din[22] ^ 
                   din[20] ^ din[19] ^ din[16] ^ din[15] ^ din[14] ^ din[12] ^ din[11] ^ 
                   din[8]  ^ din[7]  ^ din[3]  ^ cin[0]  ^ cin[3]  ^ cin[4]  ^ cin[6]  ^ 
                   cin[7]  ^ cin[9]  ^ cin[11] ^ cin[12] ^ cin[13] ^ cin[15];

  assign crc[9]  = din[30] ^ din[29] ^ din[28] ^ din[26] ^ din[24] ^ din[23] ^ din[21] ^ 
                   din[20] ^ din[17] ^ din[16] ^ din[15] ^ din[13] ^ din[12] ^ din[9]  ^ 
                   din[8]  ^ din[4]  ^ cin[0]  ^ cin[1]  ^ cin[4]  ^ cin[5]  ^ cin[7]  ^ 
                   cin[8]  ^ cin[10] ^ cin[12] ^ cin[13] ^ cin[14];

  assign crc[10] = din[31] ^ din[30] ^ din[29] ^ din[27] ^ din[25] ^ din[24] ^ din[22] ^ 
                   din[21] ^ din[18] ^ din[17] ^ din[16] ^ din[14] ^ din[13] ^ din[10] ^ 
                   din[9]  ^ din[5]  ^ cin[0]  ^ cin[1]  ^ cin[2]  ^ cin[5]  ^ cin[6]  ^ 
                   cin[8]  ^ cin[9]  ^ cin[11] ^ cin[13] ^ cin[14] ^ cin[15];

  assign crc[11] = din[31] ^ din[30] ^ din[28] ^ din[26] ^ din[25] ^ din[23] ^ din[22] ^ 
                   din[19] ^ din[18] ^ din[17] ^ din[15] ^ din[14] ^ din[11] ^ din[10] ^ 
                   din[6]  ^ cin[1]  ^ cin[2]  ^ cin[3]  ^ cin[6]  ^ cin[7]  ^ cin[9]  ^ 
                   cin[10] ^ cin[12] ^ cin[14] ^ cin[15];

  assign crc[12] = din[31] ^ din[29] ^ din[28] ^ din[24] ^ din[23] ^ din[22] ^ din[18] ^ 
                   din[16] ^ din[15] ^ din[8]  ^ din[7]  ^ din[4]  ^ din[0]  ^ cin[0]  ^ 
                   cin[2]  ^ cin[6]  ^ cin[7]  ^ cin[8]  ^ cin[12] ^ cin[13] ^ cin[15];

  assign crc[13] = din[30] ^ din[29] ^ din[25] ^ din[24] ^ din[23] ^ din[19] ^ din[17] ^ 
                   din[16] ^ din[9]  ^ din[8]  ^ din[5]  ^ din[1]  ^ cin[0]  ^ cin[1]  ^ 
                   cin[3]  ^ cin[7]  ^ cin[8]  ^ cin[9]  ^ cin[13] ^ cin[14];

  assign crc[14] = din[31] ^ din[30] ^ din[26] ^ din[25] ^ din[24] ^ din[20] ^ din[18] ^ 
                   din[17] ^ din[10] ^ din[9]  ^ din[6]  ^ din[2]  ^ cin[1]  ^ cin[2]  ^ 
                   cin[4]  ^ cin[8]  ^ cin[9]  ^ cin[10] ^ cin[14] ^ cin[15];

  assign crc[15] = din[31] ^ din[27] ^ din[26] ^ din[25] ^ din[21] ^ din[19] ^ din[18] ^ 
                   din[11] ^ din[10] ^ din[7]  ^ din[3]  ^ cin[2]  ^ cin[3]  ^ cin[5]  ^ 
                   cin[9]  ^ cin[10] ^ cin[11] ^ cin[15];
endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/phy/phy_cfg/srio_gen2_v4_1_16_phy_cfg_top.v#1 $
//----------------------------------------------------------------------
//
// PHY_CFG
// Description:
// This module contains the configuration registers for the PHY layer.
//
// It uses an AXI-Lite interface to the Configuration Fabric, and has a
// core interface for transfer of control and status information.
//
// No clock relationship between the cfg_clk and the phy_clk is
// assumed.
//
// LINK_WIDTH | PHY_CLK's relationship to gt_pcs_clk
// x4         | = gt_pcs_clk
// x2         | = gt_pcs_clk/2
// x1/trained | = gt_pcs_clk/4
//
// Hierarchy:
// PHY_TOP
//  |______PHY_CFG_TOP <-- this module
//            |______CFG_AXI (in hdl/common/)
//            |______PHY_CFG_REG
// ---------------------------------------------------------------------
`timescale 1ps/1ps
// ------------------------------------------------
// below attribute is added to supress the synthesis warnings in vivado tool 8:3332
(* DowngradeIPIdentifiedWarnings="yes" *)
// ------------------------------------------------


module srio_gen2_v4_1_16_phy_cfg_top
  #(
    parameter TCQ   = 100,
    parameter PHY_EF_PTR    = 16'h0100,   // Location of PHY  ext features {0x0100+}
    parameter LANE_EF_PTR   = 16'h0400,   // Location of Lane ext features {0x0400+}
    parameter VC_EF_PTR     = 16'h0800,   // Location of VC   ext features {0x0800+} (only if VC==1)
    parameter USER_EF_PTR   = 16'h0000,   // Location of User ext features {0x0000 or 0x0900+}
    parameter LINK_TIMEOUT  = 24'hFF_FFFF,// Link timeout ctr {0x000000-0xffffff}
    parameter PORT_TIMEOUT  = 24'hFF_FFFF,// Port timeout ctr {0x000000-0xffffff}
    parameter SW_CSR        = 0,          // SW assisted error recovery enabled {0,1}
    parameter VC            = 0,          // Highest numbered VC supported {0,1}
    parameter VC1_CT        = 1,          // Default traffic mode for VC1 (1 is CT mode) {0,1}
    parameter IS_HOST       = 1,          // Default Host value {0,1}
    parameter MASTER_EN     = 1,          // Default Master Enable value {0,1}
    parameter DISCOVERED    = 1,          // Default Discovered value {0,1}
    parameter IDLE1         = 1,          // Include IDLE1 Generator {0,1}
    parameter IDLE2         = 0,          // Include IDLE2 Generator {0,1}
    parameter MODE_XG       = 5,          // Default Line Rate {1, 2, 3, 5, 6}
    parameter GT_BYTES      = 5,          // Width of GT interface in bytes {1, 2, 4}
    parameter LINK_WIDTH    = 1)          // Number of GT lanes to use {1, 2, 4}
  (
    // {{{ Port Declarations ---------------
    // System Signals
    input             phy_clk,                // PHY interface clock
    input             phy_rst,                // Reset for PHY clock Domain
    input             gt_pcs_clk,                 // GT interface clock
    input             gt_pcs_rst,                 // Reset for GT clock domain
    input             cfg_clk,                // CFG Interface user clock
    input             cfg_rst,                // Reset for CFG clk domain

    // User Interface
    output     [23:0] PC_port_timeout,        // Timeout value user can use to detect lost packet
    output            PC_srio_host,           // Endpoint is the system host

    // LOG Interface
    output            PC_maint_only,          // LOG can only send maintenance packets
    output            PC_master_enable,       // Enable Request transactions

    // Buffer Interface
    input             BT_tx_flow_control,     // Port negotiated to tx flow control

    // OLLM TX Interface
    input      [5:0]  PT_phy_next_fm,         // Next Transmit AckID
    output     [5:0]  PC_next_fm,             // AckID to update phy_next_fm
    output     [2:0]  PC_lreq_cmd,            // Command field for Link Request
    output            PC_send_lreq,           // Register Request to send Link Request
    output            PC_load_ackids,         // Load phy_next_fm, phy_last_ack, with CFG values
    output            PC_load_nextpkt,        // Load next_rcvd_pkt with CFG value

    // OLLM RX Interface
    input      [5:0]  PR_phy_last_ack,        // Last ackID accepted by the link partner
    input      [5:0]  PR_next_rcvd_pkt,       // Next expected packet into the OLLM RX
    input      [4:0]  PR_rcvd_port_stat,      // Link partner's port status from the last received Link Response
    input      [5:0]  PR_ackid_status,        // Link partner's ackid status from the last received Link Response
    input             PR_rcvd_lresp,          // OLLM RX has received a link response
    input             PR_output_retry_stop,   // Output Retry state machine in the Output Retry Stopped State
    input             PR_output_error_stop,   // Output Error state machine in the Output Error Stopped State
    input             PR_input_retry_stop,    // Input Retry state machine in the Output Retry Stopped State
    input             PR_input_error_stop,    // Input Error state machine in the Output Error Stopped State
    input             PR_rcvd_pa_or_pna,      // Received PA or PNA
    input             PR_port_error,          // Output Error state machine in the Port Error State
    output     [5:0]  PC_next_rcvd_pkt,       // Register supplied next expected packet
    output     [5:0]  PC_last_ack,            // Register supplied last packet ack'ed value
    output     [23:0] PC_link_timeout,        // Timeout value for packet acknowledgment
    output            PC_vc_ct,               // VC in Cont. Traffic mode - turn into bus if multiple VC support added
    output            PC_vc_en,               // VC is enabled - turn into bus if multiple VC support added
    output            PC_input_maint_only,    // Only maintenance packet types are allowed
    output            PC_error_disable,       // Disable Error Checking
    output            PC_clr_port_error,      // Register supplied indication to clear port error condition

    // OPLM Interface
    input      [LINK_WIDTH*2-1:0] PP_gtrx_tap_m1_status,// tap(-1) status
    input      [LINK_WIDTH*2-1:0] PP_gtrx_tap_p1_status,// tap(+1) status
    input      [LINK_WIDTH-1:0]   PP_rx_scram_en,       // Scrambling/descrambling enabled on connected port
    input      [LINK_WIDTH-1:0]   PP_lane_sync,         // Lane sync from oplm_init
    input      [LINK_WIDTH-1:0]   PP_receiver_trained,  // Connected port lane receiver trained
    input                         PP_idle_selected,     // Indicates the IDLE sequence is selected
    input                         PP_idle2_selected,    // OPLM is in IDLE2 mode
    input      [LINK_WIDTH-1:0]   PP_idle2_rcvd,        // IDLE2 CSF received
    input                         PP_mode_1x,           // oplm_init initialized to 1x
    input                         PP_rx_lane_r,         // oplm_init initialized on lane R (valid if mode_1x asserted)
    input                         PP_port_initialized,  // Port initialized
    input      [LINK_WIDTH*4-1:0] PP_rx_lane_number,    // Lane number of connected port's lane (received in CSF)
    input      [LINK_WIDTH*3-1:0] PP_rx_port_width,     // Connected port width from IDLE2 CSF
    input      [LINK_WIDTH*4-1:0] PP_gt_decode_error,   // INVALID on GT RX (notintable or disperr)
    output     [2:0]              PC_force_lane,        // Force traindown lanes
    output                        PC_scram_disable,     // Disable scrambling
    output                        PC_port_disable,      // Port should remain in SILENT state
    output                        PC_idle2_enable,      // IDLE2 sequence is enabled

    // Configuration Fabric Interface
    input             CF_cfgp_awvalid,        // Write Address Valid
    output            PC_cfgp_awready,        // Write Address Port Ready
    input      [23:0] CF_cfgp_awaddr,         // Write Address
    input             CF_cfgp_wvalid,         // Write Data Valid
    output            PC_cfgp_wready,         // Write Data Port Ready
    input      [31:0] CF_cfgp_wdata,          // Write Data
    input      [3:0]  CF_cfgp_wstrb,          // Write Data Byte Enables
    output            PC_cfgp_bvalid,         // Write Response Valid
    input             CF_cfgp_bready,         // Write Response Fabric Ready
    input             CF_cfgp_arvalid,        // Read Address Valid
    output            PC_cfgp_arready,        // Read Address Port Ready
    input      [23:0] CF_cfgp_araddr,         // Read Address
    output            PC_cfgp_rvalid,         // Read Response Valid
    input             CF_cfgp_rready,         // Read Response Fabric Ready
    output     [31:0] PC_cfgp_rdata           // Read Data
    // }}} End Port Declarations -----------
  );

// {{{ Check Parameters ------------------
  //Catch any invalid parameter conditions
  localparam LPS_EF_SIZE  = 16'h0100;
  localparam LANE_EF_SIZE = 16'h0400;
  localparam VC_EF_SIZE   = 16'h0100;
  localparam USER_EF_SIZE = 16'h0100;

// added below macro to fix the CR# 735137
// synthesis translate_off
  initial begin
    if ((PHY_EF_PTR < 16'h0100) ||                                                            // Too small?
       (PHY_EF_PTR > (16'hffff - LPS_EF_SIZE - LANE_EF_SIZE - VC_EF_SIZE - USER_EF_SIZE)) ||  // Too big?
       (PHY_EF_PTR % LPS_EF_SIZE != 0))                                                       // Wrong boundary?
    begin
      $display("Invalid phy_ef_ptr");
      $display(PHY_EF_PTR);
      $finish; // PHY_EF_PTR is invalid
    end
    if ((LANE_EF_PTR < (PHY_EF_PTR + LPS_EF_SIZE)) ||                                         // Too small?
      (LANE_EF_PTR > (16'hffff - LANE_EF_SIZE - VC_EF_SIZE - USER_EF_SIZE)) ||               // Too big?
       (LANE_EF_PTR % LANE_EF_SIZE != 0))                                                     // Wrong boundary?
    begin
      $display("Invalid phy_ef_ptr");
      $display(LANE_EF_PTR);
      $finish; // LANE_EF_PTR is invalid
    end
    if (VC != 0) begin
      if ((VC_EF_PTR < (LANE_EF_PTR + LANE_EF_SIZE)) ||                                       // Too small?
         (VC_EF_PTR > (16'hffff - VC_EF_SIZE - USER_EF_SIZE)) ||                              // Too big?
         (VC_EF_PTR % VC_EF_SIZE != 0))                                                       // Wrong boundary?
      begin
        $finish; // VC_EF_PTR is invalid
      end
    end
    if (USER_EF_PTR > 0) begin
      if ((USER_EF_PTR < (LANE_EF_PTR + LANE_EF_SIZE + VC_EF_SIZE)) ||                        // Too small?
         (USER_EF_PTR > (16'hffff - USER_EF_SIZE)) ||                                         // Too big?
         (USER_EF_PTR % USER_EF_SIZE != 0))                                                   // Wrong boundary?
      begin
        $finish; // USER_EF_PTR is invalid
      end
    end
  end
  // }}} End Check Parameters --------------
// synthesis translate_on

  // {{{ Wire Declarations -----------------
  wire              CCA_sync_cfg_rst;         // cfg_rst sync'ed to phy_clk
  wire       [23:0] CCA_cfg_waddr;            // Write Address
  wire       [31:0] CCA_cfg_wdata;            // Write Data
  wire       [3:0]  CCA_cfg_wstrb;            // Write Data Byte Enables
  wire              CCA_sync_we;              // Synchronized write enable
  wire       [23:0] CCA_cfg_raddr;            // Read Address
  wire              CCA_sync_re;              // Synchronized Read Enable
  wire       [31:0] PCR_core_rdata;           // Read Data
  // }}} End Wire Declarations -------------

  // {{{ cfg_axi inst ----------------------
  // Instantiate the generic cfg interface, which contains the clock domain
  // crossing from cfg_clk to phy_clk, as well as the AXI-Lite interface to
  // the CFG Fabric
  srio_gen2_v4_1_16_cfg_axi
    #(
      .TCQ                       (TCQ))
    phy_cfg_axi_inst
     (.core_clk                  (phy_clk),
      .cfg_clk                   (cfg_clk),
      .cfg_rst                   (cfg_rst),
      .CF_awvalid                (CF_cfgp_awvalid),
      .CCA_awready               (PC_cfgp_awready),
      .CF_awaddr                 (CF_cfgp_awaddr),
      .CF_wvalid                 (CF_cfgp_wvalid),
      .CCA_wready                (PC_cfgp_wready),
      .CF_wdata                  (CF_cfgp_wdata),
      .CF_wstrb                  (CF_cfgp_wstrb),
      .CCA_bvalid                (PC_cfgp_bvalid),
      .CF_bready                 (CF_cfgp_bready),
      .CF_arvalid                (CF_cfgp_arvalid),
      .CCA_arready               (PC_cfgp_arready),
      .CF_araddr                 (CF_cfgp_araddr),
      .CCA_rvalid                (PC_cfgp_rvalid),
      .CF_rready                 (CF_cfgp_rready),
      .CCA_rdata                 (PC_cfgp_rdata),
      .CCA_sync_cfg_rst          (CCA_sync_cfg_rst),
      .CCA_cfg_waddr             (CCA_cfg_waddr),
      .CCA_cfg_wdata             (CCA_cfg_wdata),
      .CCA_cfg_wstrb             (CCA_cfg_wstrb),
      .CCA_sync_we               (CCA_sync_we),
      .CCA_cfg_raddr             (CCA_cfg_raddr),
      .CCA_sync_re               (CCA_sync_re),
      .CC_core_rdata             (PCR_core_rdata));
  // }}} End cfg_axi inst ------------------

  // {{{ phy_cfg_reg inst ------------------
  // Instantiate the PHY CFG register bank, containing all the CSRs for the PHY
  // layer and the interfaces to other PHY modules.
  srio_gen2_v4_1_16_phy_cfg_reg
    #(
      .TCQ                       (TCQ),
      .PHY_EF_PTR                (PHY_EF_PTR),
      .LANE_EF_PTR               (LANE_EF_PTR),
      .VC_EF_PTR                 (VC_EF_PTR),
      .USER_EF_PTR               (USER_EF_PTR),
      .LINK_TIMEOUT              (LINK_TIMEOUT),
      .PORT_TIMEOUT              (PORT_TIMEOUT),
      .SW_CSR                    (SW_CSR),
      .VC                        (VC),
      .VC1_CT                    (VC1_CT),
      .IS_HOST                   (IS_HOST),
      .MASTER_EN                 (MASTER_EN),
      .DISCOVERED                (DISCOVERED),
      .IDLE1                     (IDLE1),
      .IDLE2                     (IDLE2),
      .MODE_XG                   (MODE_XG),
      .GT_BYTES                  (GT_BYTES),
      .LINK_WIDTH                (LINK_WIDTH))
    phy_cfg_reg_inst
     (.phy_clk                   (phy_clk),
      .phy_rst                   (phy_rst),
      .gt_pcs_clk                (gt_pcs_clk),
      .gt_pcs_rst                (gt_pcs_rst),
      .CCA_sync_cfg_rst          (CCA_sync_cfg_rst),
      .PCR_port_timeout          (PC_port_timeout),
      .PCR_srio_host             (PC_srio_host),
      .PCR_maint_only            (PC_maint_only),
      .PCR_master_enable         (PC_master_enable),
      .BT_tx_flow_control        (BT_tx_flow_control),
      .PT_phy_next_fm            (PT_phy_next_fm),
      .PCR_next_fm               (PC_next_fm),
      .PCR_lreq_cmd              (PC_lreq_cmd),
      .PCR_send_lreq             (PC_send_lreq),
      .PCR_load_ackids           (PC_load_ackids),
      .PCR_load_nextpkt          (PC_load_nextpkt),
      .PR_phy_last_ack           (PR_phy_last_ack),
      .PR_next_rcvd_pkt          (PR_next_rcvd_pkt),
      .PR_rcvd_lresp             (PR_rcvd_lresp),
      .PR_ackid_status           (PR_ackid_status),
      .PR_rcvd_port_stat         (PR_rcvd_port_stat),
      .PR_output_retry_stop      (PR_output_retry_stop),
      .PR_output_error_stop      (PR_output_error_stop),
      .PR_input_retry_stop       (PR_input_retry_stop),
      .PR_input_error_stop       (PR_input_error_stop),
      .PR_rcvd_pa_or_pna         (PR_rcvd_pa_or_pna),
      .PR_port_error             (PR_port_error),
      .PCR_next_rcvd_pkt         (PC_next_rcvd_pkt),
      .PCR_last_ack              (PC_last_ack),
      .PCR_link_timeout          (PC_link_timeout),
      .PCR_vc_ct                 (PC_vc_ct),
      .PCR_vc_en                 (PC_vc_en),
      .PCR_input_maint_only      (PC_input_maint_only),
      .PCR_error_disable         (PC_error_disable),
      .PCR_clr_port_error        (PC_clr_port_error),
      .PP_gtrx_tap_m1_status     (PP_gtrx_tap_m1_status),
      .PP_gtrx_tap_p1_status     (PP_gtrx_tap_p1_status),
      .PP_rx_scram_en            (PP_rx_scram_en),
      .PP_lane_sync              (PP_lane_sync),
      .PP_receiver_trained       (PP_receiver_trained),
      .PP_idle_selected          (PP_idle_selected),
      .PP_idle2_selected         (PP_idle2_selected),
      .PP_idle2_rcvd             (PP_idle2_rcvd),
      .PP_mode_1x                (PP_mode_1x),
      .PP_rx_lane_r              (PP_rx_lane_r),
      .PP_port_initialized       (PP_port_initialized),
      .PP_rx_lane_number         (PP_rx_lane_number),
      .PP_rx_port_width          (PP_rx_port_width),
      .PP_gt_decode_error        (PP_gt_decode_error),
      .PCR_force_lane            (PC_force_lane),
      .PCR_scram_disable         (PC_scram_disable),
      .PCR_port_disable          (PC_port_disable),
      .PCR_idle2_enable          (PC_idle2_enable),
      .CCA_cfg_waddr             (CCA_cfg_waddr),
      .CCA_cfg_wdata             (CCA_cfg_wdata),
      .CCA_cfg_wstrb             (CCA_cfg_wstrb),
      .CCA_sync_we               (CCA_sync_we),
      .CCA_cfg_raddr             (CCA_cfg_raddr),
      .CCA_sync_re               (CCA_sync_re),
      .PCR_core_rdata            (PCR_core_rdata));
  // }}} End phy_cfg_reg inst --------------

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/phy/phy_cfg/srio_gen2_v4_1_16_phy_cfg_reg.v#1 $
//----------------------------------------------------------------------
//
// PHY_CFG_REG
// Description:
// This module contains the configuration registers for the PHY layer.
//
// For writes, it takes a write enable, address, data and strobe (byte
// enables) from the cfg_axi module and handles writes to writable
// registers. For reads, it takes an address and read enable, and
// returns the read data from the corresponding CSR. It also has a phy
// core interface for transfer of control and status information.
//
// No clock relationship between cfg_clk and the phy_clk is assumed.
//
// LINK_WIDTH | PHY_CLK's relationship to gt_pcs_clk
// x4         | = gt_pcs_clk*2
// x2         | = gt_pcs_clk
// x1/trained | = gt_pcs_clk/2
//
// Hierarchy:
// PHY_TOP
//    |______PHY_CFG_TOP
//              |______CFG_AXI (in hdl/common/)
//              |______PHY_CFG_REG <-- this module
// ---------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_phy_cfg_reg
  #(
    parameter TCQ   = 100,
    parameter PHY_EF_PTR    = 16'h0100,   // Location of PHY  ext features {0x0100+}
    parameter LANE_EF_PTR   = 16'h0400,   // Location of Lane ext features {0x0400+}
    parameter VC_EF_PTR     = 16'h0800,   // Location of VC   ext features {0x0800+} (only if VC==1)
    parameter USER_EF_PTR   = 16'h0000,   // Location of User ext features {0x0000 or 0x0900+}
    parameter LINK_TIMEOUT  = 24'hFF_FFFF,// Link timeout ctr {0x000000-0xffffff}
    parameter PORT_TIMEOUT  = 24'hFF_FFFF,// Port timeout ctr {0x000000-0xffffff}
    parameter SW_CSR        = 0,          // SW assisted error recovery enabled {0,1}
    parameter VC            = 0,          // Highest numbered VC supported {0,1}
    parameter VC1_CT        = 1,          // Default traffic mode for VC1 (1 is CT mode) {0,1}
    parameter IS_HOST       = 1,          // Default Host value {0,1}
    parameter MASTER_EN     = 1,          // Default Master Enable value {0,1}
    parameter DISCOVERED    = 1,          // Default Discovered value {0,1}
    parameter IDLE1         = 1,          // Include IDLE1 Generator {0,1}
    parameter IDLE2         = 0,          // Include IDLE2 Generator {0,1}
    parameter MODE_XG       = 5,          // Default Line Rate {1, 2, 3, 5, 6}
    parameter GT_BYTES      = 4,          // Width of GT interface in bytes {1, 2, 4}
    parameter LINK_WIDTH    = 1)          // Number of GT lanes to use {1, 2, 4}
  (
    // {{{ Port Declarations ---------------
    // System Signals
    input             phy_clk,                // PHY interface clock
    input             phy_rst,                // Reset for PHY clock Domain
    input             gt_pcs_clk,             // GT interface clock
    input             gt_pcs_rst,             // Reset for GT clock domain
    input             CCA_sync_cfg_rst,       // cfg_rst sync'ed to phy_clk

    // User Interface
    output reg [23:0] PCR_port_timeout = PORT_TIMEOUT,      // Timeout value user can use to detect lost packet
    output reg        PCR_srio_host = (IS_HOST == 1),       // Endpoint is the system host

    // LOG Interface
    output reg        PCR_maint_only = 1'b0,                // LOG can only send maintenance packets
    output reg        PCR_master_enable = (MASTER_EN == 1), // Enable Request transactions

    // Buffer Interface
    input             BT_tx_flow_control,                   // Port negotiated to tx flow control

    // OLLM TX Interface
    input      [5:0]  PT_phy_next_fm,                       // Next Transmit AckID
    output reg [5:0]  PCR_next_fm = 6'b0,                   // AckID to updated phy_next_fm
    output reg [2:0]  PCR_lreq_cmd = 3'b0,                  // Command field for Link Request
    output reg        PCR_send_lreq = 1'b0,                 // Register Request to send Link Request
    output reg        PCR_load_ackids = 1'b0,               // Load phy_next_fm, phy_last_ack, with CFG values
    output reg        PCR_load_nextpkt = 1'b0,              // Load next_rcvd_pkt with CFG value

    // OLLM RX Interface
    input      [5:0]  PR_phy_last_ack,                      // Last ackID accepted by the link partner
    input      [5:0]  PR_next_rcvd_pkt,                     // Next expected packet into the OLLM RX
    input             PR_rcvd_lresp,                        // OLLM RX has received a Link Response
    input      [4:0]  PR_rcvd_port_stat,                    // Link partner's port status from the Link Response
    input      [5:0]  PR_ackid_status,                      // Link partner's ackID status from the Link Response
    input             PR_output_retry_stop,                 // Output Retry fsm in the Output Retry Stopped State
    input             PR_output_error_stop,                 // Output Error fsm in the Output Error Stopped State
    input             PR_input_retry_stop,                  // Input Retry fsm in the Output Retry Stopped State
    input             PR_input_error_stop,                  // Input Error fsm in the Output Error Stopped State
    input             PR_rcvd_pa_or_pna,                    // Received PA or PNA
    input             PR_port_error,                        // Output Error state machine in the Port Error State
    output reg [5:0]  PCR_next_rcvd_pkt = 6'b0,             // Register supplied next expected packet
    output reg [5:0]  PCR_last_ack = 6'b0,                  // Register supplied last packet ack'ed value
    output reg [23:0] PCR_link_timeout = LINK_TIMEOUT,      // Timeout value for packet acknowledgment
    output reg        PCR_vc_ct =((VC == 1)&&(VC1_CT == 1)),// VC in CT mode (expand to bus if mult VC support added)
    output reg        PCR_vc_en = (VC == 1),                // VC is enabled (expand to bus if mult VC support added)
    output reg        PCR_input_maint_only = 1'b0,          // Only maintenance packet types are allowed
    output reg        PCR_error_disable = 1'b0,             // Disable Error Checking
    output reg        PCR_clr_port_error = 1'b0,            // Register supplied indication to clear port error

    // OPLM Interface
    input      [LINK_WIDTH*2-1:0] PP_gtrx_tap_m1_status,    // tap(-1) status
    input      [LINK_WIDTH*2-1:0] PP_gtrx_tap_p1_status,    // tap(+1) status
    input      [LINK_WIDTH-1:0]   PP_rx_scram_en,           // Scrambling/descrambling enabled on connected port
    input      [LINK_WIDTH-1:0]   PP_lane_sync,             // Lane sync from oplm_init
    input      [LINK_WIDTH-1:0]   PP_receiver_trained,      // Connected port lane receiver trained
    input                         PP_idle_selected,         // Indicates the IDLE sequence is selected
    input                         PP_idle2_selected,        // OPLM is in IDLE2 mode
    input      [LINK_WIDTH-1:0]   PP_idle2_rcvd,            // IDLE2 CSF received
    input                         PP_mode_1x,               // oplm_init initialized to 1x
    input                         PP_rx_lane_r,             // oplm_init initialized on lane R (valid if mode_1x asserted)
    input                         PP_port_initialized,      // Port initialized
    input      [LINK_WIDTH*4-1:0] PP_rx_lane_number,        // Lane number of connected port's lane (received in CSF)
    input      [LINK_WIDTH*3-1:0] PP_rx_port_width,         // Connected port width from IDLE2 CSF
    input      [LINK_WIDTH*4-1:0] PP_gt_decode_error,       // INVALID on GT RX (notintable or disperr)
    output reg [2:0]              PCR_force_lane    = 3'b0, // Force traindown lanes
    output reg                    PCR_scram_disable = 1'b0, // Disable scrambling
    output reg                    PCR_port_disable  = 1'b0, // Port should remain in SILENT state
    output reg                    PCR_idle2_enable  = (IDLE2 == 1),// IDLE2 sequence is enabled

    // Generic Configuration Interface
    input      [23:0] CCA_cfg_waddr,      // Write Address
    input      [31:0] CCA_cfg_wdata,      // Write Data
    input      [3:0]  CCA_cfg_wstrb,      // Write Data Byte Enables
    input             CCA_sync_we,        // Synchronized write enable
    input      [23:0] CCA_cfg_raddr,      // Read Address
    input             CCA_sync_re,        // Synchronized Read Enable
    output reg [31:0] PCR_core_rdata      // Read Data
    // }}} End Port Declarations -----------
  );

  // {{{ Localparams -----------------------
  // Parameters for the Extended Features Block IDs
  localparam LPS_EF_ID     = ((SW_CSR == 1) ? 16'h0002 : 16'h0001);   // EF_ID of LP-Serial {1, 2}
  localparam LANE_EF_ID    = 16'h000D;                                // EF_ID of LP-Serial Lane {D}
  localparam VC_EF_ID      = 16'h000A;                                // EF_ID of VC {A}

  // Parameters for CSR offsets
  // LP-Serial Extended Features Block:
  localparam [15:0] LPS_000   =  PHY_EF_PTR + 16'h0000; // Serial Register Block Header
  localparam [15:0] LPS_020   =  PHY_EF_PTR + 16'h0020; // Port Link Timeout CSR
  localparam [15:0] LPS_024   =  PHY_EF_PTR + 16'h0024; // Port Response Timeout CSR
  localparam [15:0] LPS_03C   =  PHY_EF_PTR + 16'h003c; // Port General Control CSR
  localparam [15:0] LPS_040   =  PHY_EF_PTR + 16'h0040; // Port 0 Maintenance Request CSR
  localparam [15:0] LPS_044   =  PHY_EF_PTR + 16'h0044; // Port 0 Maintenance Response CSR
  localparam [15:0] LPS_048   =  PHY_EF_PTR + 16'h0048; // Port 0 Local ackID CSR
  localparam [15:0] LPS_054   =  PHY_EF_PTR + 16'h0054; // Port 0 Control 2 CSR
  localparam [15:0] LPS_058   =  PHY_EF_PTR + 16'h0058; // Port 0 Error and Status CSR
  localparam [15:0] LPS_05C   =  PHY_EF_PTR + 16'h005C; // Port 0 Control CSR
  // LP-Serial Lane Extended Features Block:
  localparam [15:0] LANE_000  = LANE_EF_PTR + 16'h0000; // Serial Lane Register Block Header
  localparam [15:0] LANE_010  = LANE_EF_PTR + 16'h0010; // Lane 0 Status 0 CSR
  localparam [15:0] LANE_014  = LANE_EF_PTR + 16'h0014; // Lane 0 Status 1 CSR
  localparam [15:0] LANE_030  = LANE_EF_PTR + 16'h0030; // Lane 1 Status 0 CSR
  localparam [15:0] LANE_034  = LANE_EF_PTR + 16'h0034; // Lane 1 Status 1 CSR
  localparam [15:0] LANE_050  = LANE_EF_PTR + 16'h0050; // Lane 2 Status 0 CSR
  localparam [15:0] LANE_054  = LANE_EF_PTR + 16'h0054; // Lane 2 Status 1 CSR
  localparam [15:0] LANE_070  = LANE_EF_PTR + 16'h0070; // Lane 3 Status 0 CSR
  localparam [15:0] LANE_074  = LANE_EF_PTR + 16'h0074; // Lane 3 Status 1 CSR
  // Virtual Channel Extended Features Block:
  localparam [15:0] VC_000    =   VC_EF_PTR + 16'h0000; // Serial Lane Register Block Header
  localparam [15:0] VC_020    =   VC_EF_PTR + 16'h0020; // Port 0 VC CSR
  localparam [15:0] VC_024    =   VC_EF_PTR + 16'h0024; // Port 0 VC0 BW Allocation Register
  localparam [15:0] VC_028    =   VC_EF_PTR + 16'h0028; // Port 0 VC1 BW Allocation Register
  // }}} End Localparams -------------------

  // {{{ Wire Declarations -----------------
  reg           gt_pcs_rst_q;                 // registered version of gt_pcs_rst (gt_pcs_clk domain)
                                              // placeholder - not using registered version of phy_rst (phy_clk domain)
  reg           sync_cfg_rst_q;               // Registered version of CCA_sync_cfg_rst
  reg           sync_cfg_rst_ext;             // Extended cfg_rst to be used in gt_clk domain in case phy_clk > gt_clk
  reg   [7:0]   tap_m1_status;                // tap(-1) status
  reg   [7:0]   tap_p1_status;                // tap(+1) status
  reg   [3:0]   rx_scram_en;                  // scrambling/descrambling enabled on connected port
  reg   [3:0]   lane_sync;                    // lane sync from oplm_init
  reg   [3:0]   lane_sync_q;                  // registered version of lane_sync, used to detect changes in the signal
  reg   [3:0]   receiver_trained;             // connected port lane receiver trained
  reg   [11:0]  rx_port_width;                // port width from IDLE2 CSF
  reg   [3:0]   idle2_rcvd;                   // IDLE2 CSF received
  reg   [3:0]   idle2_rcvd_q;                 // registered version of idle2_rcvd, used to detect a falling edge
  wire  [3:0]   idle2_rcvd_fall;              // falling edge of idle2_rcvd (means that all CSF info is current
  reg           idle_selected;                // The core has trained to an IDLE sequence (idle2_selected is valid)
  reg           idle2_selected;               // IDLE2 operation
  reg   [15:0]  gt_decode_error;              // per lane GT decode error monitor
  reg           mode_1x;                      // oplm_init initialized to 1x
  reg           rx_lane_r;                    // oplm_init initialized to lane R
  reg           port_initialized;             // port initialized
  reg   [15:0]  rx_lane_number;               // lane number of connected port's lane (received in CSF, 4 bits/lane)
  reg           tx_flow_ctrl;                 // transmit buffer in TX flow control mode
  reg   [5:0]   phy_next_fm;                  // ackID to updated phy_next_fm
  reg   [5:0]   phy_last_ack;                 // last ackID accepted by the link partner
  wire  [5:0]   phy_last_ack_incr;            // phy_last_ack + 1
  wire  [5:0]   outstanding_ackid;            // next expected ackID for rcvd ACK control symbol (unacknowledged ackID)
  reg   [5:0]   phy_next_rcvd_pkt;            // next expected packet into the OLLM RX
  reg           output_retry_stop;            // output port in output retry-stopped state
  reg           output_error_stop;            // output port in output error-stopped state
  reg           input_retry_stop;             // input port in input retry-stopped state
  reg           input_error_stop;             // input port in input error-stopped state
  reg           port_error;                   // oplm in port error state
  reg   [2:0]   force_lane;                   // force oplm to 1x, on lane 0 or lane R
  reg           scram_disable;                // disable scrambling in oplm
  reg           port_disable;                 // force port to remain in SILENT
  reg           lane0_idle2_rcvd, lane1_idle2_rcvd, lane2_idle2_rcvd, lane3_idle2_rcvd ;  // per-lane IDLE2 indicator
  reg           lane_014_idle2_rcvd, lane_034_idle2_rcvd, lane_054_idle2_rcvd, lane_074_idle2_rcvd; // for use in CSR
  reg           idle2_enable;                 // allow IDLE2 operation (phy_clk domain)
  reg           lps_03c_discovered;           // port discovered (to user)
  reg           rcvd_lresp;                   // received link-response
  reg   [4:0]   rcvd_port_status;             // port_status from link-response
  reg   [5:0]   rcvd_ackid_status;            // ackID_status from link-response
  reg   [5:0]   ackid_status;                 // ackID status from link-response control symbol
  reg   [4:0]   link_status;                  // link status from link-response control symbol
  reg           lps_044_resp_valid;           // link-response received; status fields are valid (clr on read)
  wire  [3:0]   lps_054_baudrate;             // selected baudrate (1 - 1.25, 2 - 2.5, 3 - 3.125, 4 - 5.0, 5 - 6.25)
  reg           rcvd_pa_or_pna;               // received a packet-accepted or packet-not-accepted control symbol
  reg           lps_058_output_retried;       // output port has received a packet-retry and can not make progress
  reg           lps_058_output_retry_enc;     // output port has encountered a retry condition
  reg           lps_058_output_error_enc;     // output port has encountered a transmission error
  reg           lps_058_input_error_enc;      // input port has encountered a transmission error
  reg   [2:0]   lps_05c_init_port_width;      // initialized port width
  reg   [2:0]   port_width_ovrd_temp;         // store written port width override as it is checked for validity
  reg   [2:0]   lps_05c_port_width_ovrd;      // validated port width override
  reg           lps_05c_enum_bound;           // enumeration boundary from Port Control CSR
  reg   [3:0]   lane0_decode_error_cnt, lane1_decode_error_cnt; // Number of GT errors on this beat
  reg   [3:0]   lane2_decode_error_cnt, lane3_decode_error_cnt; // Number of GT errors on this beat
  wire  [3:0]   lane0_gt_error_cnt_d, lane1_gt_error_cnt_d;     // Cumulative GT error counters, pre-register
  wire  [3:0]   lane2_gt_error_cnt_d, lane3_gt_error_cnt_d;     // Cumulative GT error counters, pre-register
  reg   [3:0]   lane0_gt_error_cnt, lane1_gt_error_cnt;         // Cumulative GT error counters
  reg   [3:0]   lane2_gt_error_cnt, lane3_gt_error_cnt;         // Cumulative GT error counters
  reg   [3:0]   lane_sync_chg;                // lane_sync has changed
  reg   [3:0]   idle2_current;                // IDLE2 CSF information current (no errors or lane_sync state changes)
  reg   [3:0]   idle2_values_chg;             // values from the CSF have changed since Lane n Status 1 CSR was read
                // Cat of values in Lane n Status 1 CSR, and registered version of such
  wire  [14:0]  lane0_status1_csr, lane1_status1_csr, lane2_status1_csr, lane3_status1_csr;
  reg   [14:0]  lane0_status1_csr_q, lane1_status1_csr_q, lane2_status1_csr_q, lane3_status1_csr_q;
                // CSR was read
  reg           lps_044_read, lane_010_read, lane_030_read, lane_050_read, lane_070_read;
  reg           lane_014_read, lane_034_read, lane_054_read, lane_074_read;
  wire          lane_010_read_ext, lane_030_read_ext, lane_050_read_ext, lane_070_read_ext;
  wire          lane_014_read_ext, lane_034_read_ext, lane_054_read_ext, lane_074_read_ext;
  reg           lane_010_read_q, lane_030_read_q, lane_050_read_q, lane_070_read_q;
  reg           lane_014_read_q, lane_034_read_q, lane_054_read_q, lane_074_read_q;
                // CSR is being written (timing different then "CSR was read" signals)
  wire          lps_020_write, lps_024_write, lps_03c_write, lps_040_write, lps_048_write;
  wire          lps_054_write, lps_058_write, lps_05c_write, lane_014_write, lane_034_write;
  wire          lane_054_write, lane_074_write, vc_020_write;
                // Wires representing each CSR for ease of use in simulation
  wire  [31:0]  csr_lps_000, csr_lps_020, csr_lps_024, csr_lps_03c, csr_lps_040, csr_lps_044, csr_lps_048, csr_lps_054;
  wire  [31:0]  csr_lps_058, csr_lps_05c, csr_lane_000, csr_lane_010, csr_lane_014, csr_lane_030, csr_lane_034;
  wire  [31:0]  csr_lane_050, csr_lane_054, csr_lane_070, csr_lane_074, csr_vc_000, csr_vc_020, csr_vc_024, csr_vc_028;
  // }}} End Wire Declarations -------------

  // {{{ Reset Fanout Control --------------
  // Register gt_pcs_rst before use
  always @(posedge gt_pcs_clk) begin
    gt_pcs_rst_q <=  #TCQ gt_pcs_rst;
  end

  // Extend the cfg reset in case phy_clk is 2x gt_pcs_clk
  always @(posedge phy_clk) begin
    sync_cfg_rst_q   <=  #TCQ CCA_sync_cfg_rst;
    sync_cfg_rst_ext <=  #TCQ CCA_sync_cfg_rst || sync_cfg_rst_q;
  end
  // }}} End Reset Fanout Control ----------

  //   {{{ OPLM Sync -----------------------
  // Synchronize OPLM Interface (gt_pcs_clk is an integer multiple of phy_clk)

  // Register inputs in gt_pcs_clk domain, they can be used directly in phy_clk
  // domain due to clock relationship
  // These are semi-static signals
  always @(posedge gt_pcs_clk) begin
    // Unnecessary to have reset value since they're assigned from inputs on
    // every cycle
    tap_m1_status    <= #TCQ  (LINK_WIDTH == 4) ?        PP_gtrx_tap_m1_status  :
                              (LINK_WIDTH == 2) ? {4'b0, PP_gtrx_tap_m1_status} :
                              (LINK_WIDTH == 1) ? {6'b0, PP_gtrx_tap_m1_status} :
                                                   8'bx;
    tap_p1_status    <= #TCQ  (LINK_WIDTH == 4) ?        PP_gtrx_tap_p1_status  :
                              (LINK_WIDTH == 2) ? {4'b0, PP_gtrx_tap_p1_status} :
                              (LINK_WIDTH == 1) ? {6'b0, PP_gtrx_tap_p1_status} :
                                                   8'bx;
    rx_scram_en      <= #TCQ  (LINK_WIDTH == 4) ?        PP_rx_scram_en  :
                              (LINK_WIDTH == 2) ? {2'b0, PP_rx_scram_en} :
                              (LINK_WIDTH == 1) ? {3'b0, PP_rx_scram_en} :
                                                   4'bx;
    receiver_trained <= #TCQ  (LINK_WIDTH == 4) ?        PP_receiver_trained  :
                              (LINK_WIDTH == 2) ? {2'b0, PP_receiver_trained} :
                              (LINK_WIDTH == 1) ? {3'b0, PP_receiver_trained} :
                                                   4'bx;
    idle2_selected   <= #TCQ PP_idle2_selected;
    idle_selected    <= #TCQ PP_idle_selected;
    mode_1x          <= #TCQ PP_mode_1x;
    port_initialized <= #TCQ PP_port_initialized;
    rx_lane_r        <= #TCQ PP_rx_lane_r;
    rx_lane_number   <= #TCQ  (LINK_WIDTH == 4) ?         PP_rx_lane_number  :
                              (LINK_WIDTH == 2) ? {8'b0,  PP_rx_lane_number} :
                              (LINK_WIDTH == 1) ? {12'b0, PP_rx_lane_number} :
                                                   16'bx;
    rx_port_width    <= #TCQ  (LINK_WIDTH == 4) ?        PP_rx_port_width  :
                              (LINK_WIDTH == 2) ? {6'b0, PP_rx_port_width} :
                              (LINK_WIDTH == 1) ? {9'b0, PP_rx_port_width} :
                                                   12'bx;
  end

  // Same thing, but use reset value on gt_decode_error, idle2_rcvd, and
  // lane_sync to avoid X propagation
  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      gt_decode_error   <= #TCQ 16'b0;
      lane_sync         <= #TCQ 4'b0;
      lane_sync_q       <= #TCQ 4'b0;
      idle2_rcvd        <= #TCQ 4'b0;
      idle2_rcvd_q      <= #TCQ 4'b0;
    end else begin
      gt_decode_error   <= #TCQ  (LINK_WIDTH == 4) ?         PP_gt_decode_error  :
                                 (LINK_WIDTH == 2) ? {8'b0,  PP_gt_decode_error} :
                                 (LINK_WIDTH == 1) ? {12'b0, PP_gt_decode_error} :
                                                      16'bx;
      lane_sync         <= #TCQ  (LINK_WIDTH == 4) ?        PP_lane_sync  :
                                 (LINK_WIDTH == 2) ? {2'b0, PP_lane_sync} :
                                 (LINK_WIDTH == 1) ? {3'b0, PP_lane_sync} :
                                                      4'bx;
      lane_sync_q       <= #TCQ lane_sync;
      idle2_rcvd        <= #TCQ PP_idle2_rcvd;
      idle2_rcvd_q      <= #TCQ idle2_rcvd;
    end
  end

  // Register OPLM interface outputs in gt_pcs_clk domain
  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      PCR_force_lane    <= #TCQ 3'b0;
      PCR_scram_disable <= #TCQ 1'b0;
      PCR_port_disable  <= #TCQ 1'b0;
      PCR_idle2_enable  <= #TCQ (IDLE2 == 1);
    end else begin
      PCR_force_lane    <= #TCQ force_lane;
      PCR_scram_disable <= #TCQ scram_disable;
      PCR_port_disable  <= #TCQ port_disable;
      PCR_idle2_enable  <= #TCQ idle2_enable;
    end
  end
  //   }}} End OPLM Sync -------------------

  //   {{{ Other PHY modules Fanout Ctrl----
  // Outputs to core have already been registered in phy_clk domain
  // Register non-OPLM core inputs in phy_clk domain (inputs registered so that
  // phy_cfg can be located on core periphery)
  always @(posedge phy_clk) begin
    // Unnecessary to have reset value since they're assigned from inputs on
    // every cycle
    tx_flow_ctrl        <= #TCQ BT_tx_flow_control;
    phy_next_fm         <= #TCQ PT_phy_next_fm;
    phy_last_ack        <= #TCQ PR_phy_last_ack;
    phy_next_rcvd_pkt   <= #TCQ PR_next_rcvd_pkt;
    rcvd_port_status    <= #TCQ PR_rcvd_port_stat;
    rcvd_lresp          <= #TCQ PR_rcvd_lresp;
    rcvd_ackid_status   <= #TCQ PR_ackid_status;
    output_retry_stop   <= #TCQ PR_output_retry_stop;
    output_error_stop   <= #TCQ PR_output_error_stop;
    input_retry_stop    <= #TCQ PR_input_retry_stop;
    input_error_stop    <= #TCQ PR_input_error_stop;
    rcvd_pa_or_pna      <= #TCQ PR_rcvd_pa_or_pna;
    port_error          <= #TCQ PR_port_error;
  end
  //   }}} End Core Sync -------------------
  // }}} End Synchronization ---------------

  // {{{ Writable Register Bank ------------
  // A shadow register is kept for writable registers so that read and write
  // functionality can be fully separated.

  // Create signals indicating that the register is being written
  assign lps_020_write  = CCA_sync_we && (CCA_cfg_waddr[15:0] == LPS_020);
  assign lps_024_write  = CCA_sync_we && (CCA_cfg_waddr[15:0] == LPS_024);
  assign lps_03c_write  = CCA_sync_we && (CCA_cfg_waddr[15:0] == LPS_03C);
  assign lps_040_write  = CCA_sync_we && (CCA_cfg_waddr[15:0] == LPS_040);
  assign lps_048_write  = CCA_sync_we && (CCA_cfg_waddr[15:0] == LPS_048);
  assign lps_054_write  = CCA_sync_we && (CCA_cfg_waddr[15:0] == LPS_054);
  assign lps_058_write  = CCA_sync_we && (CCA_cfg_waddr[15:0] == LPS_058);
  assign lps_05c_write  = CCA_sync_we && (CCA_cfg_waddr[15:0] == LPS_05C);
  assign lane_014_write = CCA_sync_we && (CCA_cfg_waddr[15:0] == LANE_014);
  assign lane_034_write = CCA_sync_we && (CCA_cfg_waddr[15:0] == LANE_034);
  assign lane_054_write = CCA_sync_we && (CCA_cfg_waddr[15:0] == LANE_054);
  assign lane_074_write = CCA_sync_we && (CCA_cfg_waddr[15:0] == LANE_074);
  assign vc_020_write   = CCA_sync_we && (CCA_cfg_waddr[15:0] == VC_020);


  // --------------- LP-Serial Extended Features Block ------------------------
  // ----- Port Link Timeout CSR writable register(s) ----- //
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      PCR_link_timeout                <= #TCQ LINK_TIMEOUT;
    end else if (lps_020_write) begin
      if (CCA_cfg_wstrb[3])
        PCR_link_timeout[23:16]       <= #TCQ CCA_cfg_wdata[31:24];
      if (CCA_cfg_wstrb[2])
        PCR_link_timeout[15:8]        <= #TCQ CCA_cfg_wdata[23:16];
      if (CCA_cfg_wstrb[1])
        PCR_link_timeout[7:0]         <= #TCQ CCA_cfg_wdata[15:8];
    end
  end

  // ----- Port Response Timeout CSR writable register(s) ----- //
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      PCR_port_timeout                <= #TCQ PORT_TIMEOUT;
    end else if (lps_024_write) begin
      if (CCA_cfg_wstrb[3])
        PCR_port_timeout[23:16]       <= #TCQ CCA_cfg_wdata[31:24];
      if (CCA_cfg_wstrb[2])
        PCR_port_timeout[15:8]        <= #TCQ CCA_cfg_wdata[23:16];
      if (CCA_cfg_wstrb[1])
        PCR_port_timeout[7:0]         <= #TCQ CCA_cfg_wdata[15:8];
    end
  end

  // ----- Port General Control CSR writable register(s) ----- //
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      PCR_srio_host                   <= #TCQ IS_HOST;
      PCR_master_enable               <= #TCQ MASTER_EN;
      lps_03c_discovered              <= #TCQ DISCOVERED;
    end else if (lps_03c_write) begin
      if (CCA_cfg_wstrb[3]) begin
        PCR_srio_host                 <= #TCQ CCA_cfg_wdata[31];
        PCR_master_enable             <= #TCQ CCA_cfg_wdata[30];
        lps_03c_discovered            <= #TCQ CCA_cfg_wdata[29];
      end
    end
  end

  // ----- Port 0 Maintenance Request CSR writable register(s) ----- //
  //*ASSERTION*
  //(ap_send_lreq_pulse_on_write): PCR_send_lreq asserts for one cycle on write to byte 0 of Maint Req CSR
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      PCR_send_lreq                   <= #TCQ 1'b0;
    end else if (SW_CSR == 0) begin
      PCR_send_lreq                   <= #TCQ 1'b0;
    end else if (lps_040_write) begin
      if (CCA_cfg_wstrb[0]) begin
        PCR_send_lreq                 <= #TCQ 1'b1; // Pulse PCR_send_lreq high one cycle if byte 0 is written
      end
    end else begin
      PCR_send_lreq                   <= #TCQ 1'b0;
    end
  end

  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      PCR_lreq_cmd                    <= #TCQ 3'b0;
    end else if (SW_CSR == 0) begin
      PCR_lreq_cmd                    <= #TCQ 3'b0;
    end else if (lps_040_write) begin
      if (CCA_cfg_wstrb[0]) begin
        PCR_lreq_cmd                  <= #TCQ CCA_cfg_wdata[2:0]; // Update with command for LREQ
      end
    end
  end

  // ----- Port 0 Local ackID CSR writable register(s) ----- //
  //*COVERPOINT*
  //(cg_local_ackid): Group to check that Local ackIDbytes 0 and 3 are written with and without bit 31 being written
  //(cp_write_clr_outstanding_ackids): Write to Clr_outstanding_ackIDs (bit 31 = 1) in Local ackID CSR with SW_CSR = 1
  //(cp_write_inbound_ackids): Write to Inbound_ackID (byte 3) in Local ackID CSR with SW_CSR = 1
  //(cp_write_outbound_ackids): Write to Outbound_ackID (byte 0) in Local ackID CSR with SW_CSR = 1

  //*CROSS*
  //(cr_clr_ackids_and_outbound_ackids): Write to Outbound_ackID crossed with write to Clr_outstanding_ackIDs
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      PCR_next_rcvd_pkt               <= #TCQ 6'b0;
      PCR_next_fm                     <= #TCQ 6'b0;
      PCR_last_ack                    <= #TCQ 6'b0;
    end else if (SW_CSR == 0) begin
      PCR_next_rcvd_pkt               <= #TCQ 6'b0;
      PCR_next_fm                     <= #TCQ 6'b0;
      PCR_last_ack                    <= #TCQ 6'b0;
    // Ignore writes until IDLE mode trained so that ackID width is known
    end else if (lps_048_write && idle_selected) begin
      if (CCA_cfg_wstrb[3] && CCA_cfg_wdata[31]) begin
        // Clr_outstanding_ackIDs - ignore other written bits
        PCR_next_rcvd_pkt             <= #TCQ phy_next_rcvd_pkt;
        PCR_next_fm                   <= #TCQ phy_next_fm;
        PCR_last_ack                  <= #TCQ phy_next_fm - 1'b1;
      end else begin
        if (CCA_cfg_wstrb[3]) begin
          // Write to Inbound_ackID (and not Clr_outstanding_ackIDs)
          PCR_next_rcvd_pkt           <= #TCQ CCA_cfg_wdata[29:24];
        end else begin
          PCR_next_rcvd_pkt           <= #TCQ phy_next_rcvd_pkt;
        end
        if (CCA_cfg_wstrb[0]) begin
          // Write to Outbound_ackID (and not Clr_outstanding_ackIDs)
          PCR_next_fm                 <= #TCQ CCA_cfg_wdata[5:0];
          PCR_last_ack                <= #TCQ CCA_cfg_wdata[5:0] - 1'b1;
        end else begin
          PCR_next_fm                 <= #TCQ phy_next_fm;
          PCR_last_ack                <= #TCQ phy_last_ack;
        end
      end
    end
  end

  //*ASSERTION*
  //(ap_load_ackids_pulse_on_write): PCR_load_ackids high 1 cycle on write to Clr_outstanding_ackIDs or Outbound_ackID
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      PCR_load_ackids                 <= #TCQ 1'b0;
    end else if (SW_CSR == 0) begin
      PCR_load_ackids                 <= #TCQ 1'b0;
    end else if (lps_048_write && idle_selected) begin
      // PCR_load_ackids asserts one cycle if Clr_outstanding_ackIDs or Outbound_ackID is written
      if ((CCA_cfg_wstrb[3] && CCA_cfg_wdata[31]) || CCA_cfg_wstrb[0]) begin
        PCR_load_ackids               <= #TCQ 1'b1;
      end
    end else begin
      PCR_load_ackids <= #TCQ 1'b0;
    end
  end

  //*ASSERTION*
  //(ap_load_nextpkt_pulse_on_write): PCR_load_nextpkt high 1 cycle on write Inbound_ackID and !Clr_outstanding_ackIDs
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      PCR_load_nextpkt                <= #TCQ 1'b0;
    end else if (SW_CSR == 0) begin
      PCR_load_nextpkt                <= #TCQ 1'b0;
    end else if (lps_048_write && idle_selected) begin
      // PCR_load_nextpkt asserts one cycle if Inbound_ackID and is written and Clr_outstanding_ackIDs is 0
      if (CCA_cfg_wstrb[3] && !CCA_cfg_wdata[31]) begin
        PCR_load_nextpkt              <= #TCQ 1'b1;
      end
    end else begin
      PCR_load_nextpkt                <= #TCQ 1'b0;
    end
  end

  // ----- Port 0 Control 2 CSR writable register(s) ----- //
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      scram_disable                   <= #TCQ 1'b0;
    end else if (IDLE2 == 0) begin
      scram_disable                   <= #TCQ 1'b0;
    end else begin
      if (lps_054_write) begin
        if (CCA_cfg_wstrb[0]) begin
          scram_disable               <= #TCQ CCA_cfg_wdata[2];
        end
      end
    end
  end

  // ----- Port 0 Error and Status CSR writable register(s) ----- //
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      idle2_enable                    <= #TCQ (IDLE2 == 1);
    end else if (!IDLE2 || !IDLE1 || (MODE_XG > 5)) begin
      idle2_enable                    <= #TCQ (IDLE2 == 1);
    end else if (lps_058_write) begin
      if (CCA_cfg_wstrb[3]) begin
        idle2_enable                  <= #TCQ  CCA_cfg_wdata[30];
      end
    end
  end

  //*COVERPOINT*
  //(cp_clr_output_retried): Output Retried is cleared by PA or PNA
  //*ASSERTION*
  //(ap_set_clr_output_retried): Output Retried set and clear conditions do not happen together (protocol error)
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      lps_058_output_retried          <= #TCQ 1'b0;
    end else if (output_retry_stop) begin
       lps_058_output_retried         <= #TCQ 1'b1;
    end else if (rcvd_pa_or_pna) begin
       lps_058_output_retried         <= #TCQ 1'b0;
    end
  end

  //*COVERPOINT*
  //(cp_clr_output_retry_enc): Output Retry-encountered is written with 1'b1 while set
  //(cp_set_clr_output_retry_enc): Output Retry-encountered set and clr conditions happen together
  //*ASSERTION*
  //(ap_clr_output_retry_enc): lps_058_output_retry_enc is cleared when written with 1'b1
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      lps_058_output_retry_enc        <= #TCQ 1'b0;
    end else if (output_retry_stop) begin
      lps_058_output_retry_enc        <= #TCQ 1'b1;
    end else if (lps_058_write) begin
      if (CCA_cfg_wstrb[2]) begin
        if (CCA_cfg_wdata[20]) begin
          lps_058_output_retry_enc    <= #TCQ 1'b0; // Clear if written with a 1'b1
        end
      end
    end
  end

  //*COVERPOINT*
  //(cp_clr_output_error_enc): Output Error-encountered is written with 1'b1 while set
  //(cp_set_clr_output_error_enc): Output Error-encountered set and clr conditions happen together
  //*ASSERTION*
  //(ap_clr_output_error_enc): lps_058_output_error_enc is cleared when written with 1'b1
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      lps_058_output_error_enc        <= #TCQ 1'b0;
    end else if (output_error_stop) begin
      lps_058_output_error_enc        <= #TCQ 1'b1;
    end else if (lps_058_write) begin
      if (CCA_cfg_wstrb[2]) begin
        if (CCA_cfg_wdata[17]) begin
          lps_058_output_error_enc    <= #TCQ 1'b0; // Clear if written with a 1'b1
        end
      end
    end
  end

  //*COVERPOINT*
  //(cp_clr_input_error_enc): Input Error-encountered is written with 1'b1 while set
  //(cp_set_clr_input_error_enc): Input Error-encountered set and clr happen together
  //*ASSERTION*
  //(ap_clr_input_error_enc): lps_058_input_error_enc is cleared when written with 1'b1
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      lps_058_input_error_enc         <= #TCQ 1'b0;
    end else if (input_error_stop) begin
      lps_058_input_error_enc         <= #TCQ 1'b1;
    end else if (lps_058_write) begin
      if (CCA_cfg_wstrb[1]) begin
        if (CCA_cfg_wdata[9]) begin
          lps_058_input_error_enc     <= #TCQ 1'b0; // Clear if written with a 1'b1
        end
      end
    end
  end

  //*COVERPOINT*
  //(cp_clr_port_error): Port Error is written with 1'b1 while in port error state
  //*ASSERTION*
  //(ap_PCR_clr_port_error): PCR_clr_port_error is asserted for one phy_clk when written with 1'b1
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      PCR_clr_port_error              <= #TCQ 1'b0;
    end else if (lps_058_write) begin
      if (CCA_cfg_wstrb[0]) begin
        PCR_clr_port_error            <= #TCQ CCA_cfg_wdata[2]; // Assert one cycle if written with 1'b1
      end
    end else begin
      PCR_clr_port_error              <= #TCQ 1'b0;
    end
  end

  // ----- Port 0 Control CSR writable register(s) ----- //
  //*COVERPOINT*
  //(cp_unsupported_port_width_ovrd): Port Width override field written with unsupported value
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      port_width_ovrd_temp            <= #TCQ 3'b0;
      port_disable                    <= #TCQ 1'b0;
      PCR_maint_only                  <= #TCQ 1'b0;
      PCR_input_maint_only            <= #TCQ 1'b0;
      PCR_error_disable               <= #TCQ 1'b0;
      lps_05c_enum_bound              <= #TCQ 1'b0;
    end else if (lps_05c_write) begin
      if (CCA_cfg_wstrb[3])
        port_width_ovrd_temp          <= #TCQ  CCA_cfg_wdata[26:24];
      if (CCA_cfg_wstrb[2]) begin
        port_disable                  <= #TCQ  CCA_cfg_wdata[23];
        PCR_maint_only                <= #TCQ ~CCA_cfg_wdata[22];
        PCR_input_maint_only          <= #TCQ ~CCA_cfg_wdata[21];
        PCR_error_disable             <= #TCQ  CCA_cfg_wdata[20];
        lps_05c_enum_bound            <= #TCQ  CCA_cfg_wdata[17];
      end
    end
  end

  // ------------- LP-Serial Lane Extended Features Block ---------------------
  // ----- Lane 0 Status 1 CSR writable register(s) ----- //
  //*COVERAGE*
  //(cp_lane0_idle2_rcvd): lane_014_idle2_rcvd set condition occurs
  //(cp_set_clr_lane_014_idle2_rcvd): lane_014_idle2_rcvd set and clr happen together
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      lane_014_idle2_rcvd             <= #TCQ 1'b0;
    end else if (IDLE2 == 0) begin
      lane_014_idle2_rcvd             <= #TCQ 1'b0;
    end else begin
      if (lane0_idle2_rcvd) begin
        lane_014_idle2_rcvd           <= #TCQ 1'b1;
      end else if (lane_014_write) begin
        if (CCA_cfg_wstrb[3]) begin
          if (CCA_cfg_wdata[31]) // Clear if written with a 1'b1
            lane_014_idle2_rcvd       <= #TCQ 1'b0;
        end
      end
    end
  end

  // ----- Lane 1 Status 1 CSR writable register(s) ----- //
  //*COVERAGE*
  //(cp_lane1_idle2_rcvd): lane_034_idle2_rcvd set condition occurs
  //(cp_set_clr_lane_034_idle2_rcvd): lane_034_idle2_rcvd set and clr happen together
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      lane_034_idle2_rcvd             <= #TCQ 1'b0;
    end else if ((LINK_WIDTH < 2) || (IDLE2 == 0)) begin
      lane_034_idle2_rcvd             <= #TCQ 1'b0;
    end else begin
      if (lane1_idle2_rcvd) begin
        lane_034_idle2_rcvd           <= #TCQ 1'b1;
      end else if (lane_034_write) begin
        if (CCA_cfg_wstrb[3]) begin
          if (CCA_cfg_wdata[31]) // Clear if written with a 1'b1
            lane_034_idle2_rcvd       <= #TCQ 1'b0;
        end
      end
    end
  end

  // ----- Lane 2 Status 1 CSR writable register(s) ----- //
  //*COVERAGE*
  //(cp_lane2_idle2_rcvd): lane_054_idle2_rcvd set condition occurs
  //(cp_set_clr_lane_054_idle2_rcvd): lane_054_idle2_rcvd set and clr happen together
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      lane_054_idle2_rcvd             <= #TCQ 1'b0;
    end else if ((LINK_WIDTH < 4) || (IDLE2 == 0)) begin
      lane_054_idle2_rcvd             <= #TCQ 1'b0;
    end else begin
      if (lane2_idle2_rcvd) begin
        lane_054_idle2_rcvd           <= #TCQ 1'b1;
      end else if (lane_054_write) begin
        if (CCA_cfg_wstrb[3]) begin
          if (CCA_cfg_wdata[31]) // Clear if written with a 1'b1
            lane_054_idle2_rcvd       <= #TCQ 1'b0;
        end
      end
    end
  end

  // ----- Lane 3 Status 1 CSR writable register(s) ----- //
  //*COVERAGE*
  //(cp_lane3_idle2_rcvd): lane_074_idle2_rcvd set condition occurs
  //(cp_set_clr_lane_074_idle2_rcvd): lane_074_idle2_rcvd set and clr happen together
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      lane_074_idle2_rcvd             <= #TCQ 1'b0;
    end else if ((LINK_WIDTH < 4) || (IDLE2 == 0)) begin
      lane_074_idle2_rcvd             <= #TCQ 1'b0;
    end else begin
      if (lane3_idle2_rcvd) begin
        lane_074_idle2_rcvd           <= #TCQ 1'b1;
      end else if (lane_074_write) begin
        if (CCA_cfg_wstrb[3]) begin
          if (CCA_cfg_wdata[31]) // Clear if written with a 1'b1
            lane_074_idle2_rcvd       <= #TCQ 1'b0;
        end
      end
    end
  end

  // ------------ Virtual Channel Extended Features Block ---------------------
  // ----- Port 0 VC CSR writable register(s) ----- //
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      PCR_vc_ct                       <= #TCQ (VC == 1) ? VC1_CT : 1'b0;
      PCR_vc_en                       <= #TCQ (VC == 1);
    end else if (VC == 0) begin
      PCR_vc_ct                       <= #TCQ 1'b0;
      PCR_vc_en                       <= #TCQ 1'b0;
    end else if (vc_020_write) begin
      if (CCA_cfg_wstrb[2]) begin
        PCR_vc_ct                     <= #TCQ CCA_cfg_wdata[16];
      end
      if (CCA_cfg_wstrb[0]) begin
        PCR_vc_en                     <= #TCQ CCA_cfg_wdata[0];
      end
    end
  end
  // }}} End Writable Register Bank ---------

  // {{{ Gather Information For Read -------
  // Create signals needed for registers

  //   {{{ phy_clk domain signals ----------
  // Calculate phy_last_ack + 1 for use in several registers
  assign phy_last_ack_incr = phy_last_ack + 1'b1;

  // Mask off upper bit of phy_last_ack_incr in IDLE1 operation
  assign outstanding_ackid = {(idle2_selected && phy_last_ack_incr[5]),phy_last_ack_incr[4:0]};

  // Port 0 Control CSR - Port Width Support field
  assign lps_054_baudrate = MODE_XG == 1 ? 4'b0001 : // 1.25 GBaud
                            MODE_XG == 2 ? 4'b0010 : // 2.5 GBaud
                            MODE_XG == 3 ? 4'b0011 : // 3.125 GBaud
                            MODE_XG == 5 ? 4'b0100 : // 5.0 GBaud
                            MODE_XG == 6 ? 4'b0101 : // 6.25 GBaud
                                           4'b0000 ; // no rate selected - spec indicates this is reset value,
                                                     // but because of parameter checking, we should never see this

  // Port 0 Link Maintenance CSR response_valid field
  // Clear on read, set when LRESP is received
  //*COVERPOINT*
  //(cp_rcvd_lresp_and_read): Receive LRESP while LPS_044 being read
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      lps_044_resp_valid       <= #TCQ 1'b0;
    end else if (SW_CSR == 1) begin
      if (rcvd_lresp) begin
        lps_044_resp_valid     <= #TCQ 1'b1;
      end else if (lps_044_read) begin
        lps_044_resp_valid     <= #TCQ 1'b0;
      end
    end
  end

  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      link_status   <= #TCQ 5'b0;
      ackid_status  <= #TCQ 6'b0;
    end else if (SW_CSR == 0) begin
      link_status   <= #TCQ 5'b0;
      ackid_status  <= #TCQ 6'b0;
    end else if (rcvd_lresp) begin
      link_status   <= #TCQ rcvd_port_status;
      ackid_status  <= #TCQ rcvd_ackid_status;
    end
  end


  // Port 0 Control CSR port width override field
  // Allow writing of only supported values based on LINK_WIDTH
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      lps_05c_port_width_ovrd <= #TCQ 3'b0;
    end else begin
      case (LINK_WIDTH)
        1: begin
          case (port_width_ovrd_temp)
            3'b000, 3'b010 :                  lps_05c_port_width_ovrd  <= #TCQ port_width_ovrd_temp;
            default :                         lps_05c_port_width_ovrd  <= #TCQ lps_05c_port_width_ovrd;
          endcase
        end
        2: begin
          case (port_width_ovrd_temp)
            3'b000, 3'b010, 3'b011, 3'b101 :  lps_05c_port_width_ovrd  <= #TCQ port_width_ovrd_temp;
            default :                         lps_05c_port_width_ovrd  <= #TCQ lps_05c_port_width_ovrd;
          endcase
        end
        4: begin
          case (port_width_ovrd_temp)
            3'b000, 3'b010, 3'b011, 3'b110 :  lps_05c_port_width_ovrd  <= #TCQ port_width_ovrd_temp;
            default :                         lps_05c_port_width_ovrd  <= #TCQ lps_05c_port_width_ovrd;
          endcase
        end
      endcase
    end
  end

  // Drive force lane based on port width override
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      force_lane      <= #TCQ 3'b0;
    end else begin
      force_lane  <= #TCQ lps_05c_port_width_ovrd;
    end
  end
  //   }}} phy_clk domain signals ----------

  //   {{{ gt_pcs_clk domain signals -----------
  // Port 0 Control CSR initialized port width field
  always @(posedge gt_pcs_clk) begin
    // Do not use a reset since the spec allows for it to be 'implementation dependent'
    lps_05c_init_port_width  <= #TCQ      (mode_1x &&  rx_lane_r)  ? 3'b001 : // Single-lane port, lane R
                    ((LINK_WIDTH == 1) || (mode_1x && !rx_lane_r)) ? 3'b000 : // Single-lane port
                    ((LINK_WIDTH == 4) && !mode_1x)                ? 3'b010 : // Four-lane port
                    ((LINK_WIDTH == 2) && !mode_1x)                ? 3'b011 : // Two-lane port
                                                                     3'bxxx ; // Undefined
  end

  // Lane n Status 0 CSRs 8B/10B decoding errors
  // Saturating 4-bit binary counter in gt_pcs_clk domain, inc for each byte with an error

  always @(posedge gt_pcs_clk) begin
//    if (sync_cfg_rst_ext) begin
    if (CCA_sync_cfg_rst) begin
      lane0_decode_error_cnt <= #TCQ 4'b0;
      lane1_decode_error_cnt <= #TCQ 4'b0;
      lane2_decode_error_cnt <= #TCQ 4'b0;
      lane3_decode_error_cnt <= #TCQ 4'b0;
    end else begin
      lane0_decode_error_cnt <= #TCQ  gt_decode_error[0] +
                                      (gt_decode_error[1] && GT_BYTES >1) +
                                      (gt_decode_error[2] && GT_BYTES >2) +
                                      (gt_decode_error[3] && GT_BYTES >3) ;
      lane1_decode_error_cnt <= #TCQ  gt_decode_error[GT_BYTES*1+0] +
                                      (gt_decode_error[GT_BYTES*1+1] && GT_BYTES >1) +
                                      (gt_decode_error[GT_BYTES*1+2] && GT_BYTES >2) +
                                      (gt_decode_error[GT_BYTES*1+3] && GT_BYTES >3) ;
      lane2_decode_error_cnt <= #TCQ  gt_decode_error[GT_BYTES*2+0] +
                                      (gt_decode_error[GT_BYTES*2+1] && GT_BYTES >1) +
                                      (gt_decode_error[GT_BYTES*2+2] && GT_BYTES >2) +
                                      (gt_decode_error[GT_BYTES*2+3] && GT_BYTES >3) ;
      lane3_decode_error_cnt <= #TCQ  gt_decode_error[GT_BYTES*3+0] +
                                      (gt_decode_error[GT_BYTES*3+1] && GT_BYTES >1) +
                                      (gt_decode_error[GT_BYTES*3+2] && GT_BYTES >2) +
                                      (gt_decode_error[GT_BYTES*3+3] && GT_BYTES >3) ;
    end
  end

  assign lane0_gt_error_cnt_d = lane0_decode_error_cnt + lane0_gt_error_cnt;
  assign lane1_gt_error_cnt_d = lane1_decode_error_cnt + lane1_gt_error_cnt;
  assign lane2_gt_error_cnt_d = lane2_decode_error_cnt + lane2_gt_error_cnt;
  assign lane3_gt_error_cnt_d = lane3_decode_error_cnt + lane3_gt_error_cnt;

  // Lane 0
  //*COVERPOINT*
  //(cg_gterr_ctr0): Lane 0 GT counter values
  //(cp_gt_decode_err0): Lane 0 GT decode error(s) detected
  //*CROSS*
  //(cr_gterr_full_inc0): GT decode error detected after counter saturates
  //*ASSERTION*
  //(ap_gterr_ctr0_overflow): lane0_gt_error ctr does not overflow
  always @(posedge gt_pcs_clk) begin
//    if (sync_cfg_rst_ext) begin
    if (CCA_sync_cfg_rst) begin
      lane0_gt_error_cnt            <= #TCQ 4'b0;
    end else begin
      if (lane_010_read_ext) begin                  // Clr on read (possible to miss up to 8 gt errors during read -
        lane0_gt_error_cnt          <= #TCQ 4'b0;   // lane_010_read_ext asserts one cycle after read for two phy_clks)
      end else begin
        if (lane0_gt_error_cnt[3] && !lane0_gt_error_cnt_d[3]) begin
          lane0_gt_error_cnt      <= #TCQ 4'b1111;  // Counter saturates at 4'b1111
        end else begin
          lane0_gt_error_cnt      <= #TCQ lane0_gt_error_cnt_d;
        end
      end
    end
  end
  // Lane 1
  //*COVERPOINT*
  //(cg_gterr_ctr1): Lane 1 GT counter values
  //(cp_gt_decode_err1): Lane 1 GT decode error(s) detected
  //*CROSS*
  //(cr_gterr_full_inc1): GT decode error detected after counter saturates
  //*ASSERTION*
  //(ap_gterr_ctr1_overflow): lane1_gt_error ctr does not overflow
  always @(posedge gt_pcs_clk) begin
//    if (sync_cfg_rst_ext) begin
    if (CCA_sync_cfg_rst) begin
      lane1_gt_error_cnt            <= #TCQ 4'b0;
    end else begin
      if (lane_030_read_ext) begin                  // Clr on read (possible to miss up to 8 gt errors during read -
        lane1_gt_error_cnt          <= #TCQ 4'b0;   // lane_030_read_ext asserts one cycle after read for two phy_clks)
      end else begin
        if (lane1_gt_error_cnt[3] && !lane1_gt_error_cnt_d[3]) begin
          lane1_gt_error_cnt      <= #TCQ 4'b1111;  // Counter saturates at 4'b1111
        end else begin
          lane1_gt_error_cnt      <= #TCQ lane1_gt_error_cnt_d;
        end
      end
    end
  end
  // Lane 2
  //*COVERPOINT*
  //(cg_gterr_ctr2): Lane 2 GT counter values
  //(cp_gt_decode_err2): Lane 2 GT decode error(s) detected
  //*CROSS*
  //(cr_gterr_full_inc2): GT decode error detected after counter saturates
  //*ASSERTION*
  //(ap_gterr_ctr2_overflow): lane2_gt_error ctr does not overflow
  always @(posedge gt_pcs_clk) begin
//    if (sync_cfg_rst_ext) begin
    if (CCA_sync_cfg_rst) begin
      lane2_gt_error_cnt            <= #TCQ 4'b0;
    end else begin
      if (lane_050_read_ext) begin                  // Clr on read (possible to miss up to 8 gt errors during read -
        lane2_gt_error_cnt          <= #TCQ 4'b0;   // lane_050_read_ext asserts one cycle after read for two phy_clks)
      end else begin
        if (lane2_gt_error_cnt[3] && !lane2_gt_error_cnt_d[3]) begin
          lane2_gt_error_cnt      <= #TCQ 4'b1111;  // Counter saturates at 4'b1111
        end else begin
          lane2_gt_error_cnt      <= #TCQ lane2_gt_error_cnt_d;
        end
      end
    end
  end

  // Lane 3
  //*COVERPOINT*
  //(cg_gterr_ctr3): Lane 3 GT counter values
  //(cp_gt_decode_err3): Lane 3 GT decode error(s) detected
  //*CROSS*
  //(cr_gterr_full_inc3): GT decode error detected after counter saturates
  //*ASSERTION*
  //(ap_gterr_ctr3_overflow): lane3_gt_error ctr does not overflow
  always @(posedge gt_pcs_clk) begin
//    if (sync_cfg_rst_ext) begin
    if (CCA_sync_cfg_rst) begin
      lane3_gt_error_cnt            <= #TCQ 4'b0;
    end else begin
      if (lane_070_read_ext) begin                  // Clr on read (possible to miss up to 8 gt errors during read -
        lane3_gt_error_cnt          <= #TCQ 4'b0;   // lane_070_read_ext asserts one cycle after read for two phy_clks)
      end else begin
        if (lane3_gt_error_cnt[3] && !lane3_gt_error_cnt_d[3]) begin
          lane3_gt_error_cnt      <= #TCQ 4'b1111;  // Counter saturates at 4'b1111
        end else begin
          lane3_gt_error_cnt      <= #TCQ lane3_gt_error_cnt_d;
        end
      end
    end
  end

  // Lane n Status 0 CSR's Lane_sync state change field
  // Looks for a change in lane_sync from OPLM, operates in gt_pcs_clk domain
  // The change in lane_sync takes precedence over the write-to-clear, to make
  // sure that no state changes are missed from the SW's perspective.
  //*COVERPOINT*
  //(cp_lane0_sync_chg_and_read): lane_sync for lane 0 changed while Lane 0 Status CSR was read (set & clr together)
  //(cp_lane1_sync_chg_and_read): lane_sync for lane 1 changed while Lane 0 Status CSR was read (set & clr together)
  //(cp_lane2_sync_chg_and_read): lane_sync for lane 2 changed while Lane 0 Status CSR was read (set & clr together)
  //(cp_lane3_sync_chg_and_read): lane_sync for lane 3 changed while Lane 0 Status CSR was read (set & clr together)
  always @(posedge gt_pcs_clk) begin
//    if (sync_cfg_rst_ext) begin
    if (CCA_sync_cfg_rst) begin
      lane_sync_chg          <= #TCQ 4'b0;
    end else begin
      // Lane 0
      if (lane_sync_q[0] != lane_sync[0]) begin
        lane_sync_chg[0]     <= #TCQ 1'b1;
      end else if (lane_010_read_ext) begin // clear on read; phy_clk domain signal - ok b/c of clock relationship
        lane_sync_chg[0]     <= #TCQ 1'b0;
      end
      // Lane 1
      if (lane_sync_q[1] != lane_sync[1]) begin
        lane_sync_chg[1]     <= #TCQ 1'b1;
      end else if (lane_030_read_ext) begin // clear on read; phy_clk domain signal - ok b/c of clock relationship
        lane_sync_chg[1]     <= #TCQ 1'b0;
      end
      // Lane 2
      if (lane_sync_q[2] != lane_sync[2]) begin
        lane_sync_chg[2]     <= #TCQ 1'b1;
      end else if (lane_050_read_ext) begin // clear on read; phy_clk domain signal - ok b/c of clock relationship
        lane_sync_chg[2]     <= #TCQ 1'b0;
      end
      // Lane 3
      if (lane_sync_q[3] != lane_sync[3]) begin
        lane_sync_chg[3]     <= #TCQ 1'b1;
      end else if (lane_070_read_ext) begin // clear on read; phy_clk domain signal - ok b/c of clock relationship
        lane_sync_chg[3]     <= #TCQ 1'b0;
      end
    end
  end

  // Check for falling edge of idle2_rcvd
  assign idle2_rcvd_fall = ~idle2_rcvd & idle2_rcvd_q;

  // Assign per-lane idle2_rcvd based on current port width and active lane(s)
  always @(*)
    case(LINK_WIDTH)
      1: begin
        lane0_idle2_rcvd = idle2_rcvd_fall[0];
        lane1_idle2_rcvd = 1'b0;
        lane2_idle2_rcvd = 1'b0;
        lane3_idle2_rcvd = 1'b0;
      end
      2: begin
        lane0_idle2_rcvd = ((mode_1x &&  rx_lane_r) ? 1'b0 : idle2_rcvd_fall[0]);
        lane1_idle2_rcvd = ((mode_1x && !rx_lane_r) ? 1'b0 : idle2_rcvd_fall[1]);
        lane2_idle2_rcvd = 1'b0;
        lane3_idle2_rcvd = 1'b0;
      end
      4: begin
        lane0_idle2_rcvd = ((mode_1x &&  rx_lane_r) ? 1'b0 : idle2_rcvd_fall[0]);
        lane1_idle2_rcvd = ( mode_1x                ? 1'b0 : idle2_rcvd_fall[1]);
        lane2_idle2_rcvd = ((mode_1x && !rx_lane_r) ? 1'b0 : idle2_rcvd_fall[2]);
        lane3_idle2_rcvd = ( mode_1x                ? 1'b0 : idle2_rcvd_fall[3]);
      end
      default: begin
        lane0_idle2_rcvd = 1'b0;
        lane1_idle2_rcvd = 1'b0;
        lane2_idle2_rcvd = 1'b0;
        lane3_idle2_rcvd = 1'b0;
      end
    endcase

  // Lane n Status 1 CSR's IDLE2 information current field
  // Set when IDLE2 is received and clears if lane_sync goes to '0', operates in gt_pcs_clk domain
  //*COVERPOINT*
  //(cp_not_lane0_sync_and_idle2_rcvd): IDLE2 received while lane 0 out of sync
  //(cp_not_lane1_sync_and_idle2_rcvd): IDLE2 received while lane 1 out of sync
  //(cp_not_lane2_sync_and_idle2_rcvd): IDLE2 received while lane 2 out of sync
  //(cp_not_lane3_sync_and_idle2_rcvd): IDLE2 received while lane 3 out of sync
  always @(posedge gt_pcs_clk) begin
//    if (sync_cfg_rst_ext) begin
    if (CCA_sync_cfg_rst) begin
      idle2_current           <= #TCQ 4'b0;
    end else begin
      // Lane 0
      if (!lane_sync[0]) begin
        idle2_current[0]      <= #TCQ 1'b0;
      end else if (lane0_idle2_rcvd) begin
        idle2_current[0]      <= #TCQ 1'b1;
      end
      // Lane 1
      if (!lane_sync[1]) begin
        idle2_current[1]      <= #TCQ 1'b0;
      end else if (lane1_idle2_rcvd) begin
        idle2_current[1]      <= #TCQ 1'b1;
      end
      // Lane 2
      if (!lane_sync[2]) begin
        idle2_current[2]      <= #TCQ 1'b0;
      end else if (lane2_idle2_rcvd) begin
        idle2_current[2]      <= #TCQ 1'b1;
      end
      // Lane 3
      if (!lane_sync[3]) begin
        idle2_current[3]      <= #TCQ 1'b0;
      end else if (lane3_idle2_rcvd) begin
        idle2_current[3]      <= #TCQ 1'b1;
      end
    end
  end

  // Lane n Status 1 CSRs Values changed field
  // Set if any bits in the CSR change, cleared when read

  //*ASSERTION*
  //(ap_lane0_idle2_chg_missed): No IDLE2 value changes missed on lane 0
  //(ap_lane1_idle2_chg_missed): No IDLE2 value changes missed on lane 1
  //(ap_lane2_idle2_chg_missed): No IDLE2 value changes missed on lane 2
  //(ap_lane3_idle2_chg_missed): No IDLE2 value changes missed on lane 3

  assign lane0_status1_csr = {lane_014_idle2_rcvd, idle2_current[0], receiver_trained[0],
                              rx_port_width[2:0], rx_lane_number[3:0], tap_m1_status[1:0],
                              tap_p1_status[1:0], rx_scram_en[0]};
  assign lane1_status1_csr = {lane_034_idle2_rcvd, idle2_current[1], receiver_trained[1],
                              rx_port_width[5:3], rx_lane_number[7:4], tap_m1_status[3:2],
                              tap_p1_status[3:2], rx_scram_en[1]};
  assign lane2_status1_csr = {lane_054_idle2_rcvd, idle2_current[2], receiver_trained[2],
                              rx_port_width[8:6], rx_lane_number[11:8], tap_m1_status[5:4],
                              tap_p1_status[5:4], rx_scram_en[2]};
  assign lane3_status1_csr = {lane_074_idle2_rcvd, idle2_current[3], receiver_trained[3],
                              rx_port_width[11:9], rx_lane_number[15:12], tap_m1_status[7:6],
                              tap_p1_status[7:6], rx_scram_en[3]};

  //*COVERPOINT*
  //(cp_lane0_idle2_chg_and_read): Lane 0 IDLE2 values change while being read
  //(cp_lane1_idle2_chg_and_read): Lane 1 IDLE2 values change while being read
  //(cp_lane2_idle2_chg_and_read): Lane 2 IDLE2 values change while being read
  //(cp_lane3_idle2_chg_and_read): Lane 3 IDLE2 values change while being read

  always @(posedge gt_pcs_clk) begin
//    if (sync_cfg_rst_ext) begin
    if (CCA_sync_cfg_rst) begin
      idle2_values_chg            <= #TCQ 4'hF; // spec'ed reset value to all ones (Rev 2.1 Table 6-22)

    // No reset needed on lanen_status1_csr_q signals since assigned immediately
    end else begin
      lane0_status1_csr_q         <= #TCQ lane0_status1_csr;
      lane1_status1_csr_q         <= #TCQ lane1_status1_csr;
      lane2_status1_csr_q         <= #TCQ lane2_status1_csr;
      lane3_status1_csr_q         <= #TCQ lane3_status1_csr;
      // Lane 0
      if (lane0_status1_csr != lane0_status1_csr_q) begin
        idle2_values_chg[0]      <= #TCQ 1'b1;
      end else if (lane_014_read_ext) begin // clear on read
        idle2_values_chg[0]      <= #TCQ 1'b0;
      end
      // Lane 1
      if (lane1_status1_csr != lane1_status1_csr_q) begin
        idle2_values_chg[1]      <= #TCQ 1'b1;
      end else if (lane_034_read_ext) begin // clear on read
        idle2_values_chg[1]      <= #TCQ 1'b0;
      end
      // Lane 2
      if (lane2_status1_csr != lane2_status1_csr_q) begin
        idle2_values_chg[2]      <= #TCQ 1'b1;
      end else if (lane_054_read_ext) begin // clear on read
        idle2_values_chg[2]      <= #TCQ 1'b0;
      end
      // Lane 3
      if (lane3_status1_csr != lane3_status1_csr_q) begin
        idle2_values_chg[3]      <= #TCQ 1'b1;
      end else if (lane_074_read_ext) begin // clear on read
        idle2_values_chg[3]      <= #TCQ 1'b0;
      end
    end
  end

  //   }}} gt_pcs_clk domain signals -----------
  // }}} End Gather Information For Read ---

  // {{{ Read Data Assembly ----------------
  // Form read data based on address
  // Bit ordering mirrors RapidIO Spec (e.g. spec bit 0 -> phy_cfg bit 31)
  // Note that some inputs are in the phy_clk domain, some in the gt_pcs_clk domain
  // Since gt_pcs_clk is an integer multiple of phy_clk, it is acceptable to sample
  // the signals directly in the phy_clk domain

  // Create wires for each CSR for easy simulation viewing.
  // ----------------- LP-Serial Extended Features Block --------------------------
                                                    // core  (spec)   Description
                                                    // ----------------------------
  // LP-Serial Register Block Header
  assign csr_lps_000 =  {LANE_EF_PTR[15:0],         // 31:16  (0:15)  Ptr to next EF
                         LPS_EF_ID[15:0]};          // 15:0   (16:31) LP-Serial EF_ID

  // Port Link Timeout CSR
  assign csr_lps_020 =  {PCR_link_timeout,          // 31:8   (0:23)  Link Timeout Value
                         8'b0};                     // 7:0    (24:31) Reserved

  // Port Response Timeout CSR
  assign csr_lps_024 =  {PCR_port_timeout,          // 31:8   (0:23)  Port Timeout Value
                         8'b0};                     // 7:0    (24:31) Reserved

  // Port General Control CSR
  assign csr_lps_03c =  {PCR_srio_host,             // 31     (0)     Host
                         PCR_master_enable,         // 30     (1)     Master Enable
                         lps_03c_discovered,        // 29     (2)     Discovered
                         29'b0};                    // 28:0   (3:31)  Reserved

  // Port 0 Link Maintenance Request CSR
  assign csr_lps_040 =  (SW_CSR == 0) ? 32'b0 :     //                Return 0's if unimplemented
                        {29'b0,                     // 31:3   (0:28)  Reserved
                         PCR_lreq_cmd};             // 2:0    (29:31) Link Request Command

  // Port 0 Link Maintenance Response CSR
  assign csr_lps_044 =  (SW_CSR == 0) ? 32'b0 :     //                Return 0's if unimplemented
                        {lps_044_resp_valid,        // 31     (0)     Lresp status valid
                         20'b0,                     // 30:11  (1:20)  Reserved
                         ackid_status,              // 10:5   (21:26) ackID_status
                         link_status};              // 4:0    (27:31) link_status

  // Port 0 Local ackID Status CSR
  assign csr_lps_048 =  (SW_CSR == 0) ? 32'b0 :     //                Return 0's if unimplemented
                        {2'b0,                      // 31:30  (0:1)   Clr_outstanding_ackIDs, Reserved
                         phy_next_rcvd_pkt,         // 29:24  (2:7)   Inbound_ackID
                         10'b0,                     // 23:14  (8:17)  Reserved
                         outstanding_ackid,         // 13:8   (18:23) Outstanding_ackID
                         2'b0,                      // 7:6    (24:25) Reserved
                         phy_next_fm};              // 5:0    (26:31) Outbound_ackID

  // Port 0 Control 2 CSR
  assign csr_lps_054 =  {lps_054_baudrate,          // 31:28  (0:3)   Selected Baudrate
                         2'b0,                      // 27:26  (4:5)   Reserved
                         (MODE_XG == 1),            // 25     (6)     1.25 GBaud Support
                         (MODE_XG == 1),            // 24     (7)     1.25 GBaud Enable
                         (MODE_XG == 2),            // 23     (8)     2.5 GBaud Support
                         (MODE_XG == 2),            // 22     (9)     2.5 GBaud Enable
                         (MODE_XG == 3),            // 21     (10)    3.125 GBaud Support
                         (MODE_XG == 3),            // 20     (11)    3.125 GBaud Enable
                         (MODE_XG == 5),            // 19     (12)    5.0 GBaud Support
                         (MODE_XG == 5),            // 18     (13)    5.0 GBaud Enable
                         (MODE_XG == 6),            // 17     (14)    6.25 GBaud Support
                         (MODE_XG == 6),            // 16     (15)    6.25 GBaud Enable
                         13'b0,                     // 15:3   (16:28) Reserved
                         scram_disable,             // 2      (29)    Data scrambling disable
                         2'b0};                     // 1:0    (30:31) Reserved

  // Port 0 Error and Status CSR
  assign csr_lps_058 =  {(IDLE2 == 1),              // 31     (0)     Idle Sequence 2 support
                         idle2_enable,              // 30     (1)     Idle Sequence 2 Enable
                         idle2_selected,            // 29     (2)     Idle Sequence
                         1'b0,                      // 28     (3)     Reserved
                         tx_flow_ctrl,              // 27     (4)     Flow Control Mode
                         6'b0,                      // 26:21  (5:10)  Reserved
                         lps_058_output_retry_enc,  // 20     (11)    Output Retry-encountered
                         lps_058_output_retried,    // 19     (12)    Output Retried
                         output_retry_stop,         // 18     (13)    Output Retry-stopped
                         lps_058_output_error_enc,  // 17     (14)    Output Error-encountered
                         output_error_stop,         // 16     (15)    Output Error-stopped
                         5'b0,                      // 15:11  (16:20) Reserved
                         input_retry_stop,          // 10     (21)    Input Retry-stopped
                         lps_058_input_error_enc,   // 9      (22)    Input Error-encountered
                         input_error_stop,          // 8      (23)    Input Error-stopped
                         5'b0,                      // 7:3    (24:28) Reserved, Port-write Pending, Port Unavailable
                         port_error,                // 2      (29)    Port Error
                         port_initialized,          // 1      (30)    Port OK
                         ~port_initialized};        // 0      (31)    Port Uninitialized

  // Port 0 Control CSR
  assign csr_lps_05c =  {(LINK_WIDTH == 2),         // 31     (0)     Port Width Support bit 0
                         (LINK_WIDTH == 4),         // 30     (1)     Port Width Support bit 1
                         lps_05c_init_port_width,   // 29:27  (2:4)   Initialized Port Width
                         lps_05c_port_width_ovrd,   // 26:24  (5:7)   Port Width Override
                         port_disable,              // 23     (8)     Port Disable
                         !PCR_maint_only,           // 22     (9)     Output Port Enable
                         !PCR_input_maint_only,     // 21     (10)    Input Port Enable
                         PCR_error_disable,         // 20     (11)    Error Checking Disable
                         1'b1,                      // 19     (12)    Multicast-event Participant
                         1'b0,                      // 18     (13)    Reserved
                         lps_05c_enum_bound,        // 17     (14)    Enumeration Boundary
                         16'b0,                     // 16:1   (15:30) Rsvd, Extended Port Width Support/Override
                         1'b1};                     // 0      (31)    Port Type (serial port)

  // --------------- LP-Serial Lane Extended Features Block -----------------------
                                                    // core  (spec)   Description
                                                    // ----------------------------
  // LP-Serial Lane Register Block Header
  assign csr_lane_000 = {((VC == 0) ? 
                         USER_EF_PTR[15:0] :        // 31:16  (0:15)  Ptr to next EF (VC if enabled, else user EF)
                         VC_EF_PTR[15:0]),          // 31:16  (0:15)  Ptr to next EF (VC if enabled, else user EF)
                         LANE_EF_ID[15:0]};         // 15:0   (16:31) LP-Serial Lane EF_ID

  // Lane 0 Status 0 CSR
  assign csr_lane_010 = {8'b0,                      // 31:24  (0:7)   Port Number
                        4'b0000,                    // 23:20  (8:11)  Lane Number
                        5'b0,                       // 19:15  (12:16) TX type/mode, RX type, RX input inverted
                        lane_sync[0],               // 14     (17)    Receiver trained
                        lane_sync[0],               // 13     (18)    Receiver lane sync
                        lane_sync[0],               // 12     (19)    Receiver lane ready
                        lane0_gt_error_cnt,         // 11:8   (20:23) 8B/10B decoding errors
                        lane_sync_chg[0],           // 7      (24)    Lane_sync state change
                        lane_sync_chg[0],           // 6      (25)    Rcvr_trained state change
                        2'b0,                       // 5:4    (26:27) Reserved
                        (IDLE2 == 1),               // 3      (28)    Status 1 CSR Implemented
                        3'b0};                      // 2:0    (29:31) Status 2-7 CSRs Implemented

  // Lane 0 Status 1 CSR
  assign csr_lane_014 = (IDLE2 == 0) ? 32'b0 :      //                Return 0's if unimplemented
                        {lane_014_idle2_rcvd,       // 31     (0)     IDLE2 received
                         idle2_current[0],          // 30     (1)     IDLE2 information current
                         idle2_values_chg[0],       // 29     (2)     Values Changed
                         1'b0,                      // 28     (3)     Implementation defined
                         receiver_trained[0],       // 27     (4)     Connected port lane receiver trained
                         rx_port_width[2:0],        // 26:24  (5:7)   Received port width
                         rx_lane_number[3:0],       // 23:20  (8:11)  Lane number in connected port
                         tap_m1_status[1:0],        // 19:18  (12:13) Connected port tx emphasis Tap (-1) status
                         tap_p1_status[1:0],        // 17:16  (14:15) Connected port tx emphasis Tap (+1) status
                         rx_scram_en[0],            // 15     (16)    Connected port scrambling/descrambling enabled
                         15'b0};                    // 14:0   (17:31) Reserved

  // Lane 1 Status 0 CSR
  assign csr_lane_030 = (LINK_WIDTH < 2) ? 32'b0 :  //                Return 0's if unimplemented
                        {8'b0,                      // 31:24  (0:7)   Port Number
                         4'b0001,                   // 23:20  (8:11)  Lane Number
                         5'b0,                      // 19:15  (12:16) TX type/mode, RX type, RX input inverted
                         lane_sync[1],              // 14     (17)    Receiver trained
                         lane_sync[1],              // 13     (18)    Receiver lane sync
                         lane_sync[1],              // 12     (019)   Receiver lane ready
                         lane1_gt_error_cnt,        // 11:8   (20:23) 8B/10B decoding errors
                         lane_sync_chg[1],          // 7      (24)    Lane_sync state change
                         lane_sync_chg[1],          // 6      (25)    Rcvr_trained state change
                         2'b0,                      // 5:4    (26:27) Reserved
                         (IDLE2 == 1),              // 3      (28)    Status 1 CSR Implemented
                         3'b0};                     // 2:0    (29:31) Status 2-7 CSRs Implemented

  // Lane 1 Status 1 CSR
  assign csr_lane_034 = (IDLE2 == 0) ? 32'b0 :      //                Return 0's if unimplemented
                        (LINK_WIDTH < 2) ? 32'b0 :  //                Return 0's if unimplemented
                        {lane_034_idle2_rcvd,       // 31     (0)     IDLE2 received
                         idle2_current[1],          // 30     (1)     IDLE2 information current
                         idle2_values_chg[1],       // 29     (2)     Values Changed
                         1'b0,                      // 28     (3)     Implementation defined
                         receiver_trained[1],       // 27     (4)     Connected port lane receiver trained
                         rx_port_width[5:3],        // 26:24  (5:7)   Received port width
                         rx_lane_number[7:4],       // 23:20  (8:11)  Lane number in connected port
                         tap_m1_status[3:2],        // 19:18  (12:13) Connected port tx emphasis Tap (-1) status
                         tap_p1_status[3:2],        // 17:16  (14:15) Connected port tx emphasis Tap (+1) status
                         rx_scram_en[1],            // 15     (16)    Connected port scrambling/descrambling enabled
                         15'b0};                    // 14:0   (17:31) Reserved

  // Lane 2 Status 0 CSR
  assign csr_lane_050 = (LINK_WIDTH < 4) ? 32'b0 :  //                Return 0's if unimplemented
                        {8'b0,                      // 31:24  (0:7)   Port Number
                         4'b0010,                   // 23:20  (8:11)  Lane Number
                         5'b0,                      // 19:15  (12:16) TX type/mode, RX type, RX input inverted
                         lane_sync[2],              // 14     (17)    Receiver trained
                         lane_sync[2],              // 13     (18)    Receiver lane sync
                         lane_sync[2],              // 12     (19)    Receiver lane ready
                         lane2_gt_error_cnt,        // 11:8   (20:23) 8B/10B decoding errors
                         lane_sync_chg[2],          // 7      (24)    Lane_sync state change
                         lane_sync_chg[2],          // 6      (25)    Rcvr_trained state change
                         2'b0,                      // 5:4    (26:27) Reserved
                         (IDLE2 == 1),              // 3      (28)    Status 1 CSR Implemented
                         3'b0};                     // 2:0    (29:31) Status 2-7 CSRs Implemented

  // Lane 2 Status 1 CSR
  assign csr_lane_054 = (IDLE2 == 0) ? 32'b0 :      //                Return 0's if unimplemented
                        (LINK_WIDTH < 4) ? 32'b0 :  //                Return 0's if unimplemented
                        {lane_054_idle2_rcvd,       // 31     (0)     IDLE2 received
                         idle2_current[2],          // 30     (1)     IDLE2 information current
                         idle2_values_chg[2],       // 29     (2)     Values Changed
                         1'b0,                      // 28     (3)     Implementation defined
                         receiver_trained[2],       // 27     (4)     Connected port lane receiver trained
                         rx_port_width[8:6],        // 26:24  (5:7)   Received port width
                         rx_lane_number[11:8],      // 23:20  (8:11)  Lane number in connected port
                         tap_m1_status[5:4],        // 19:18  (12:13) Connected port tx emphasis Tap (-1) status
                         tap_p1_status[5:4],        // 17:16  (14:15) Connected port tx emphasis Tap (+1) status
                         rx_scram_en[2],            // 15     (16)    Connected port scrambling/descrambling enabled
                         15'b0};                    // 14:0   (17:31) Reserved

  // Lane 3 Status 0 CSR
  assign csr_lane_070 = (LINK_WIDTH < 4) ? 32'b0 :  //                Return 0's if unimplemented
                        {8'b0,                      // 31:24  (0:7)   Port Number
                         4'b0011,                   // 23:20  (8:11)  Lane Number
                         5'b0,                      // 19:15  (12:16) TX type/mode, RX type, RX input inverted
                         lane_sync[3],              // 14     (17)    Receiver trained
                         lane_sync[3],              // 13     (18)    Receiver lane sync
                         lane_sync[3],              // 12     (19)    Receiver lane ready
                         lane3_gt_error_cnt,        // 11:8   (20:23) 8B/10B decoding errors
                         lane_sync_chg[3],          // 7      (24)    Lane_sync state change
                         lane_sync_chg[3],          // 6      (25)    Rcvr_trained state change
                         2'b0,                      // 5:4    (26:27) Reserved
                         (IDLE2 == 1),              // 3      (28)    Status 1 CSR Implemented
                         3'b0};                     // 2:0    (29:31) Status 2-7 CSRs Implemented

  // Lane 3 Status 1 CSR
  assign csr_lane_074 = (IDLE2 == 0) ? 32'b0 :      //                Return 0's if unimplemented
                        (LINK_WIDTH < 4) ? 32'b0 :  //                Return 0's if unimplemented
                        {lane_074_idle2_rcvd,       // 31     (0)     IDLE2 received
                         idle2_current[3],          // 30     (1)     IDLE2 information current
                         idle2_values_chg[3],       // 29     (2)     Values Changed
                         1'b0,                      // 28     (3)     Implementation defined
                         receiver_trained[3],       // 27     (4)     Connected port lane receiver trained
                         rx_port_width[11:9],       // 26:24  (5:7)   Received port width
                         rx_lane_number[15:12],     // 23:20  (8:11)  Lane number in connected port
                         tap_m1_status[7:6],        // 19:18  (12:13) Connected port tx emphasis Tap (-1) status
                         tap_p1_status[7:6],        // 17:16  (14:15) Connected port tx emphasis Tap (+1) status
                         rx_scram_en[3],            // 15     (16)    Connected port scrambling/descrambling enabled
                         15'b0};                    // 14:0   (17:31) Reserved

  // -------------- Virtual Channel Extended Features Block -----------------------
  // Accesses to VC Extended Features Block should retun 0's unless
  // VC is set.
                                                    // core  (spec)   Description
                                                    // ----------------------------
  // VC Register Block Header
  assign csr_vc_000   = (VC == 0) ? 32'b0 :         //                Return 0's if unimplemented
                        {USER_EF_PTR[15:0],         // 31:16  (0:15)  Ptr to next EF
                         VC_EF_ID[15:0]};           // 15:0   (16:31) Virtual Channel EF_ID

  // Port 0 VC CSR
  assign csr_vc_020   = (VC == 0) ? 32'b0 :         //                Return 0's if unimplemented
                        {8'b0,                      // 31:24  (0:7)   VC Refresh Interval
                         7'b0, PCR_vc_ct,           // 23:16  (8:15)  CT Mode
                         8'b0000_0001,              // 15:8   (16:23) VCs Support
                         7'b0, PCR_vc_en};          // 7:0    (24:31) VCs Enable

  // Port 0 VC0 BW Allocation Register
  assign csr_vc_024   = (VC == 0) ? 32'b0 :         //                Return 0's if unimplemented
                         32'b0;                     // 31:0   (0:31)  VC0 BW Allocation Reg

  // Port 0 VC 5, VC 1 BW Allocation Register
  assign csr_vc_028   = (VC == 0) ? 32'b0 :         //                Return 0's if unimplemented
                        {16'b0,                     // 31:16  (0:15)  Reserved (VC 5 is not supported)
                         16'hFF00};                 // 15:0   (16:31) BW Allocation for VC 1

  //*COVERAGE*
  //(cp_lps_000_rd_b4_wr): Cover that each byte of lps_000 was read before it was written
  //(cp_lps_000_rd_aftr_wr): Cover that each byte of lps_000 was read after it was written
  //(cp_lps_020_rd_b4_wr): Cover that each byte of lps_020 was read before it was written
  //(cp_lps_020_rd_aftr_wr): Cover that each byte of lps_020 was read after it was written
  //(cp_lps_020_3_rst_val_chk): Cover that LINK_TIMEOUT is non-default and lps_020 byte 3 was rd_b4_wr
  //(cp_lps_020_2_rst_val_chk): Cover that LINK_TIMEOUT is non-default and lps_020 byte 2 was rd_b4_wr
  //(cp_lps_020_1_rst_val_chk): Cover that LINK_TIMEOUT is non-default and lps_020 byte 1 was rd_b4_wr
  //(cp_lps_024_rd_b4_wr): Cover that each byte of lps_024 was read before it was written
  //(cp_lps_024_rd_aftr_wr): Cover that each byte of lps_024 was read after it was written
  //(cp_lps_024_3_rst_val_chk): Cover that PORT_TIMEOUT is non-default and lps_024 byte 3 was rd_b4_wr
  //(cp_lps_024_2_rst_val_chk): Cover that PORT_TIMEOUT is non-default and lps_024 byte 2 was rd_b4_wr
  //(cp_lps_024_1_rst_val_chk): Cover that PORT_TIMEOUT is non-default and lps_024 byte 1 was rd_b4_wr
  //(cp_lps_03c_rd_b4_wr): Cover that each byte of lps_03c was read before it was written
  //(cp_lps_03c_rd_aftr_wr): Cover that each byte of lps_03c was read after it was written
  //(cp_lps_03c_bit31_rst_val_chk): Cover that IS_HOST is non-default and lps_03c bit 31 was rd_b4_wr
  //(cp_lps_03c_bit30_rst_val_chk): Cover that MASTER_EN is non-default and lps_03c bit 30 was rd_b4_wr
  //(cp_lps_03c_bit29_rst_val_chk): Cover that DISCOVERED is non-default and lps_03c bit 29 was rd_b4_wr
  //(cp_lps_040_rd_b4_wr): Cover that each byte of lps_040 was read before it was written
  //(cp_lps_040_rd_aftr_wr): Cover that each byte of lps_040 was read after it was written
  //(cp_lps_044_rd_b4_wr): Cover that each byte of lps_044 was read before it was written
  //(cp_lps_044_rd_aftr_wr): Cover that each byte of lps_044 was read after it was written
  //(cp_lps_048_rd_b4_wr): Cover that each byte of lps_048 was read before it was written
  //(cp_lps_048_rd_aftr_wr): Cover that each byte of lps_048 was read after it was written
  //(cp_lps_054_rd_b4_wr): Cover that each byte of lps_054 was read before it was written
  //(cp_lps_054_rd_aftr_wr): Cover that each byte of lps_054 was read after it was written
  //(cp_lps_058_rd_b4_wr): Cover that each byte of lps_058 was read before it was written
  //(cp_lps_058_rd_aftr_wr): Cover that each byte of lps_058 was read after it was written
  //(cp_lps_058_bit30_rst_val_chk): Cover that IDLE2 is non-default and lps_058 bit 30 was rd_b4_wr
  //(cp_lps_05c_rd_b4_wr): Cover that each byte of lps_05c was read before it was written
  //(cp_lps_05c_rd_aftr_wr): Cover that each byte of lps_05c was read after it was written
  //(cp_lane_000_rd_b4_wr): Cover that each byte of lane_000 was read before it was written
  //(cp_lane_000_rd_aftr_wr): Cover that each byte of lane_000 was read after it was written
  //(cp_lane_010_rd_b4_wr): Cover that each byte of lane_010 was read before it was written
  //(cp_lane_010_rd_aftr_wr): Cover that each byte of lane_010 was read after it was written
  //(cp_lane_014_rd_b4_wr): Cover that each byte of lane_014 was read before it was written
  //(cp_lane_014_rd_aftr_wr): Cover that each byte of lane_014 was read after it was written
  //(cp_rst_lane_014_idle2_rcvd): lane_014_idle2_rcvd is reset by writing 1'b1
  //(cp_lane_030_rd_b4_wr): Cover that each byte of lane_030 was read before it was written
  //(cp_lane_030_rd_aftr_wr): Cover that each byte of lane_030 was read after it was written
  //(cp_lane_034_rd_b4_wr): Cover that each byte of lane_034 was read before it was written
  //(cp_lane_034_rd_aftr_wr): Cover that each byte of lane_034 was read after it was written
  //(cp_rst_lane_034_idle2_rcvd): lane_034_idle2_rcvd is reset by writing 1'b1
  //(cp_lane_050_rd_b4_wr): Cover that each byte of lane_050 was read before it was written
  //(cp_lane_050_rd_aftr_wr): Cover that each byte of lane_050 was read after it was written
  //(cp_lane_054_rd_b4_wr): Cover that each byte of lane_054 was read before it was written
  //(cp_lane_054_rd_aftr_wr): Cover that each byte of lane_054 was read after it was written
  //(cp_rst_lane_054_idle2_rcvd): lane_054_idle2_rcvd is reset by writing 1'b1
  //(cp_lane_070_rd_b4_wr): Cover that each byte of lane_070 was read before it was written
  //(cp_lane_070_rd_aftr_wr): Cover that each byte of lane_070 was read after it was written
  //(cp_lane_074_rd_b4_wr): Cover that each byte of lane_074 was read before it was written
  //(cp_lane_074_rd_aftr_wr): Cover that each byte of lane_074 was read after it was written
  //(cp_rst_lane_074_idle2_rcvd): lane_074_idle2_rcvd is reset by writing 1'b1
  //(cp_vc_000_rd_b4_wr): Cover that each byte of vc_000 was read before it was written
  //(cp_vc_000_rd_aftr_wr): Cover that each byte of vc_000 was read after it was written
  //(cp_vc_020_rd_b4_wr): Cover that each byte of vc_020 was read before it was written
  //(cp_vc_020_rd_aftr_wr): Cover that each byte of vc_020 was read after it was written
  //(cp_vc_020_bit16_rst_val_chk): Cover that VC and VC1_CT are non-default and vc_020 bit 16 was rd_b4_wr
  //(cp_vc_020_bit0_rst_val_chk): Cover that VC is non-default and vc_020 bit 0 was rd_b4_wr
  //(cp_vc_024_rd_b4_wr): Cover that each byte of vc_024 was read before it was written
  //(cp_vc_024_rd_aftr_wr): Cover that each byte of vc_024 was read after it was written
  //(cp_vc_028_rd_b4_wr): Cover that each byte of vc_028 was read before it was written
  //(cp_vc_028_rd_aftr_wr): Cover that each byte of vc_028 was read after it was written

  // Register read data when address is safe
  // No reset needed since data is not sampled until valid
  always @(posedge phy_clk) begin
    if (CCA_sync_re) begin
      case (CCA_cfg_raddr[15:0])
        LPS_000    : PCR_core_rdata <= #TCQ csr_lps_000;
        LPS_020    : PCR_core_rdata <= #TCQ csr_lps_020;
        LPS_024    : PCR_core_rdata <= #TCQ csr_lps_024;
        LPS_03C    : PCR_core_rdata <= #TCQ csr_lps_03c;
        LPS_040    : PCR_core_rdata <= #TCQ csr_lps_040;
        LPS_044    : PCR_core_rdata <= #TCQ csr_lps_044;
        LPS_048    : PCR_core_rdata <= #TCQ csr_lps_048;
        LPS_054    : PCR_core_rdata <= #TCQ csr_lps_054;
        LPS_058    : PCR_core_rdata <= #TCQ csr_lps_058;
        LPS_05C    : PCR_core_rdata <= #TCQ csr_lps_05c;
        LANE_000   : PCR_core_rdata <= #TCQ csr_lane_000;
        LANE_010   : PCR_core_rdata <= #TCQ csr_lane_010;
        LANE_014   : PCR_core_rdata <= #TCQ csr_lane_014;
        LANE_030   : PCR_core_rdata <= #TCQ csr_lane_030;
        LANE_034   : PCR_core_rdata <= #TCQ csr_lane_034;
        LANE_050   : PCR_core_rdata <= #TCQ csr_lane_050;
        LANE_054   : PCR_core_rdata <= #TCQ csr_lane_054;
        LANE_070   : PCR_core_rdata <= #TCQ csr_lane_070;
        LANE_074   : PCR_core_rdata <= #TCQ csr_lane_074;
        VC_000     : PCR_core_rdata <= #TCQ csr_vc_000;
        VC_020     : PCR_core_rdata <= #TCQ csr_vc_020;
        VC_024     : PCR_core_rdata <= #TCQ csr_vc_024;
        VC_028     : PCR_core_rdata <= #TCQ csr_vc_028;
        // Return data of all 0's if read to unimplemented space
        default    : PCR_core_rdata <= #TCQ 32'b0;
      endcase
    end
  end

  // Create signals to indicate register was read - used for clearing on read
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      lps_044_read  <= #TCQ 1'b0;
      lane_010_read <= #TCQ 1'b0;
      lane_014_read <= #TCQ 1'b0;
      lane_030_read <= #TCQ 1'b0;
      lane_034_read <= #TCQ 1'b0;
      lane_050_read <= #TCQ 1'b0;
      lane_054_read <= #TCQ 1'b0;
      lane_070_read <= #TCQ 1'b0;
      lane_074_read <= #TCQ 1'b0;
    end else begin
      lps_044_read  <= #TCQ CCA_sync_re && (CCA_cfg_raddr[15:0] == LPS_044);
      lane_010_read <= #TCQ CCA_sync_re && (CCA_cfg_raddr[15:0] == LANE_010);
      lane_014_read <= #TCQ CCA_sync_re && (CCA_cfg_raddr[15:0] == LANE_014);
      lane_030_read <= #TCQ CCA_sync_re && (CCA_cfg_raddr[15:0] == LANE_030);
      lane_034_read <= #TCQ CCA_sync_re && (CCA_cfg_raddr[15:0] == LANE_034);
      lane_050_read <= #TCQ CCA_sync_re && (CCA_cfg_raddr[15:0] == LANE_050);
      lane_054_read <= #TCQ CCA_sync_re && (CCA_cfg_raddr[15:0] == LANE_054);
      lane_070_read <= #TCQ CCA_sync_re && (CCA_cfg_raddr[15:0] == LANE_070);
      lane_074_read <= #TCQ CCA_sync_re && (CCA_cfg_raddr[15:0] == LANE_074);
    end
  end

  // Register read signals that will be used in the gt_pcs_clk domain so that they
  // can be extended in case phy_clk is faster than gt_pcs_clk
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      lane_010_read_q   <= #TCQ 1'b0;
      lane_014_read_q   <= #TCQ 1'b0;
      lane_030_read_q   <= #TCQ 1'b0;
      lane_034_read_q   <= #TCQ 1'b0;
      lane_050_read_q   <= #TCQ 1'b0;
      lane_054_read_q   <= #TCQ 1'b0;
      lane_070_read_q   <= #TCQ 1'b0;
      lane_074_read_q   <= #TCQ 1'b0;
    end else begin
      lane_010_read_q   <= #TCQ lane_010_read;
      lane_014_read_q   <= #TCQ lane_014_read;
      lane_030_read_q   <= #TCQ lane_030_read;
      lane_034_read_q   <= #TCQ lane_034_read;
      lane_050_read_q   <= #TCQ lane_050_read;
      lane_054_read_q   <= #TCQ lane_054_read;
      lane_070_read_q   <= #TCQ lane_070_read;
      lane_074_read_q   <= #TCQ lane_074_read;
    end
  end

  // Extend read signals for use in the gt_pcs_clk domain
  assign lane_010_read_ext = ((LINK_WIDTH == 4) && !mode_1x && lane_010_read_q) || lane_010_read;
  assign lane_014_read_ext = ((LINK_WIDTH == 4) && !mode_1x && lane_014_read_q) || lane_014_read;
  assign lane_030_read_ext = ((LINK_WIDTH == 4) && !mode_1x && lane_030_read_q) || lane_030_read;
  assign lane_034_read_ext = ((LINK_WIDTH == 4) && !mode_1x && lane_034_read_q) || lane_034_read;
  assign lane_050_read_ext = ((LINK_WIDTH == 4) && !mode_1x && lane_050_read_q) || lane_050_read;
  assign lane_054_read_ext = ((LINK_WIDTH == 4) && !mode_1x && lane_054_read_q) || lane_054_read;
  assign lane_070_read_ext = ((LINK_WIDTH == 4) && !mode_1x && lane_070_read_q) || lane_070_read;
  assign lane_074_read_ext = ((LINK_WIDTH == 4) && !mode_1x && lane_074_read_q) || lane_074_read;

  //*COVERAGE*
  //(cg_port_error_and_status_rd): Group to check that the error bits are read as 1's and 0's.
  //(cp_output_retry_enc): Cover that Output Retry-encountered was a 1 and 0 on a read
  //(cp_output_error_enc): Cover that Output Error-encountered was a 1 and 0 on a read
  //(cp_input_error_enc): Cover that Input Error-encountered was a 1 and 0 on a read

  // }}} End Read Data Assembly ------------


endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/phy/oplm/srio_gen2_v4_1_16_oplm_gtregisters.v#1 $
//----------------------------------------------------------------------
//
// OPLM_LFSR
// Description:
// This module simply registers all the inputs used from the GTs. This is 
// done in order to improve timing through the tools.  If the GT_REG 
// parameter is not set, this is bypassed.
//
// Hierarchy:
// PHY_TOP
//    |___OPLM_TOP
//            |___OPLM_GTREGISTERS <-- this module
// ---------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_oplm_gtregisters #(
    parameter TCQ           = 100,
    parameter LINK_WIDTH    = 1,                      // {1, 2, 4}
    parameter GT_BYTES      = 4,                      // GT Interface Width
    parameter DATA_WIDTH    = LINK_WIDTH*GT_BYTES*8,  // Data width
    parameter CHARIS_WIDTH  = LINK_WIDTH*GT_BYTES,    // Charisk bus width
    parameter GT_REG        = 1)                      // Indicates to register the GT inputs first
  (
    // {{{ port declarations ---------------
    // System Signals
    input                           gt_pcs_clk,      //GT Clock
    input                           gt_pcs_rst_q,    //GT reset

    //GT inputs
    input       [DATA_WIDTH-1:0]    GT_gtrx_data,           //Receive Data
    input       [CHARIS_WIDTH-1:0]  GT_gtrx_charisk,        //Character is K
    input       [CHARIS_WIDTH-1:0]  GT_gtrx_chariscomma,    //Character is Comma
    input       [CHARIS_WIDTH-1:0]  GT_gtrx_disperr,        //Disperity Error
    input       [CHARIS_WIDTH-1:0]  GT_gtrx_notintable,     //Not in Table
    input       [LINK_WIDTH-1:0]    GT_gtrx_chanisaligned,  //Channel is Aligned
    input                           GT_gtrx_reset_req,      //RX Buffer Error
    input       [LINK_WIDTH-1:0]    GT_gtrx_reset_done,     //RX Buffer Resets done
    
    //Registered Outputs
    (* shreg_extract = "no" *)
    output reg  [DATA_WIDTH-1:0]    PPG_gtrx_data,          //Receive Data
    (* shreg_extract = "no" *)
    output reg  [CHARIS_WIDTH-1:0]  PPG_gtrx_chariskchar,   //Character is K
    (* shreg_extract = "no" *)
    output reg  [CHARIS_WIDTH-1:0]  PPG_gtrx_charisa,       //Character is /A/
    (* shreg_extract = "no" *)
    output reg  [CHARIS_WIDTH-1:0]  PPG_gtrx_charisk,       //Character is /K/    
    (* shreg_extract = "no" *)
    output reg  [CHARIS_WIDTH-1:0]  PPG_gtrx_charisr,       //Character is /R/   
    (* shreg_extract = "no" *)
    output reg  [CHARIS_WIDTH-1:0]  PPG_gtrx_charism,       //Character is /M/
    (* shreg_extract = "no" *)
    output reg  [CHARIS_WIDTH-1:0]  PPG_gtrx_charispd,      //Character is /PD/
    (* shreg_extract = "no" *)
    output reg  [CHARIS_WIDTH-1:0]  PPG_gtrx_charissc,      //Character is /SC/
    (* shreg_extract = "no" *)
    output reg  [CHARIS_WIDTH-1:0]  PPG_gtrx_chariscomma,   //Character is Comma
    (* shreg_extract = "no" *)
    output reg  [CHARIS_WIDTH-1:0]  PPG_gtrx_invalid,       //Disperity Error
    (* shreg_extract = "no" *)
    output reg  [LINK_WIDTH-1:0]    PPG_gtrx_chanisaligned, //Channel is Aligned

    (* shreg_extract = "no" *)
    output reg                      PPG_gtrx_reset_req,     //RX Buffer Error 
    (* shreg_extract = "no" *)
    output reg  [LINK_WIDTH-1:0]    PPG_gtrx_reset_done     //RX Buffer Resets done
    // }}} end port declarations -----------
  );

  // Local parameter to simplify the gt interface with the data paths for 
  // character detection
  localparam A_CHAR  = 8'hFB;
  localparam K_CHAR  = 8'hBC; 
  localparam R_CHAR  = 8'hFD;
  localparam M_CHAR  = 8'h3C;
  localparam PD_CHAR = 8'h7C;
  localparam SC_CHAR = 8'h1C;

  (* shreg_extract = "no" *)
  reg  [DATA_WIDTH-1:0]       PPG_gtrx_data_d;
  (* shreg_extract = "no" *)
  reg  [CHARIS_WIDTH-1:0]     PPG_gtrx_chariskchar_d;   
  (* shreg_extract = "no" *)
  reg  [CHARIS_WIDTH-1:0]     PPG_gtrx_chariscomma_d;
  (* shreg_extract = "no" *)
  reg  [CHARIS_WIDTH-1:0]     PPG_gtrx_invalid_d;
  (* shreg_extract = "no" *)
  reg  [LINK_WIDTH-1:0]       PPG_gtrx_chanisaligned_d;
  (* shreg_extract = "no" *)
  reg                         PPG_gtrx_reset_req_d;
  (* shreg_extract = "no" *)
  reg  [LINK_WIDTH-1:0]       PPG_gtrx_reset_done_d;

  genvar ii;
  genvar jj;

  //Register the outputs if the GT_REG parameter is set
  generate if (GT_REG) begin: gtreg_gen
    // First registers the GT inputs for timing
    always @(posedge gt_pcs_clk) begin
      // need a reset on these to keep the core in sync with the testbench
      if (gt_pcs_rst_q) begin
        PPG_gtrx_data_d          <= #TCQ 0;
        PPG_gtrx_chariskchar_d   <= #TCQ 0;
        PPG_gtrx_chariscomma_d   <= #TCQ 0;
        PPG_gtrx_invalid_d       <= #TCQ 0;
        PPG_gtrx_chanisaligned_d <= #TCQ 0;
        PPG_gtrx_reset_req_d     <= #TCQ 0;
        PPG_gtrx_reset_done_d    <= #TCQ 0;
      end else begin
        PPG_gtrx_data_d          <= #TCQ GT_gtrx_data;
        PPG_gtrx_chariskchar_d   <= #TCQ GT_gtrx_charisk;
        PPG_gtrx_chariscomma_d   <= #TCQ GT_gtrx_chariscomma;
        PPG_gtrx_invalid_d       <= #TCQ GT_gtrx_disperr | GT_gtrx_notintable;
        PPG_gtrx_chanisaligned_d <= #TCQ GT_gtrx_chanisaligned;
        PPG_gtrx_reset_req_d     <= #TCQ GT_gtrx_reset_req;
        PPG_gtrx_reset_done_d    <= #TCQ GT_gtrx_reset_done;
      end
    end

    always @(posedge gt_pcs_clk) begin
      // need a reset on these to keep the core in sync with the testbench
      if (gt_pcs_rst_q) begin
        PPG_gtrx_data            <= #TCQ 0;
        PPG_gtrx_chariskchar     <= #TCQ 0;
        PPG_gtrx_chariscomma     <= #TCQ 0;
        PPG_gtrx_invalid         <= #TCQ 0;
        PPG_gtrx_chanisaligned   <= #TCQ 0;
        PPG_gtrx_reset_req       <= #TCQ 0;
        PPG_gtrx_reset_done      <= #TCQ 0;
      end else begin
        PPG_gtrx_data            <= #TCQ PPG_gtrx_data_d;
        PPG_gtrx_chariskchar     <= #TCQ PPG_gtrx_chariskchar_d;
        PPG_gtrx_chariscomma     <= #TCQ PPG_gtrx_chariscomma_d & ~PPG_gtrx_invalid_d;
        PPG_gtrx_invalid         <= #TCQ PPG_gtrx_invalid_d;
        PPG_gtrx_chanisaligned   <= #TCQ PPG_gtrx_chanisaligned_d;
        PPG_gtrx_reset_req       <= #TCQ PPG_gtrx_reset_req_d;
        PPG_gtrx_reset_done      <= #TCQ PPG_gtrx_reset_done_d;
      end
    end
    
    // Determine what characters are before passed to the init and rx modules
    // for better timing
    for (ii=0; ii < LINK_WIDTH; ii=ii+1) begin : charisx_gen
      wire [GT_BYTES-1:0] is_a;
      wire [GT_BYTES-1:0] is_k;
      wire [GT_BYTES-1:0] is_r;
      wire [GT_BYTES-1:0] is_m;
      wire [GT_BYTES-1:0] is_pd;
      wire [GT_BYTES-1:0] is_sc;

      for (jj=0; jj < GT_BYTES; jj=jj+1) begin: charisx_gtbytes_gen
        assign is_a[jj] = (PPG_gtrx_chariskchar_d[(ii*GT_BYTES)+jj] & ~PPG_gtrx_invalid_d[(ii*GT_BYTES)+jj]) &&
                          (PPG_gtrx_data_d[((ii*GT_BYTES*8)+(jj*8))+:8] == A_CHAR);

        assign is_k[jj] = (PPG_gtrx_chariskchar_d[(ii*GT_BYTES)+jj] & ~PPG_gtrx_invalid_d[(ii*GT_BYTES)+jj]) &&
                          (PPG_gtrx_data_d[((ii*GT_BYTES*8)+(jj*8))+:8] == K_CHAR);

        assign is_r[jj] = (PPG_gtrx_chariskchar_d[(ii*GT_BYTES)+jj] & ~PPG_gtrx_invalid_d[(ii*GT_BYTES)+jj]) &&
                          (PPG_gtrx_data_d[((ii*GT_BYTES*8)+(jj*8))+:8] == R_CHAR);

        assign is_m[jj] = (PPG_gtrx_chariskchar_d[(ii*GT_BYTES)+jj] & ~PPG_gtrx_invalid_d[(ii*GT_BYTES)+jj]) &&
                          (PPG_gtrx_data_d[((ii*GT_BYTES*8)+(jj*8))+:8] == M_CHAR);

        assign is_pd[jj] = (PPG_gtrx_chariskchar_d[(ii*GT_BYTES)+jj] & ~PPG_gtrx_invalid_d[(ii*GT_BYTES)+jj]) &&
                           (PPG_gtrx_data_d[((ii*GT_BYTES*8)+(jj*8))+:8] == PD_CHAR);

        assign is_sc[jj] = (PPG_gtrx_chariskchar_d[(ii*GT_BYTES)+jj] & ~PPG_gtrx_invalid_d[(ii*GT_BYTES)+jj]) &&
                           (PPG_gtrx_data_d[((ii*GT_BYTES*8)+(jj*8))+:8] == SC_CHAR);

        always @(posedge gt_pcs_clk) begin
          // need a reset on these to keep the core in sync with the testbench
          if (gt_pcs_rst_q) begin
            PPG_gtrx_charisa[ii*GT_BYTES+jj]   <= #TCQ 0;
            PPG_gtrx_charisk[ii*GT_BYTES+jj]   <= #TCQ 0;
            PPG_gtrx_charisr[ii*GT_BYTES+jj]   <= #TCQ 0;
            PPG_gtrx_charism[ii*GT_BYTES+jj]   <= #TCQ 0;
            PPG_gtrx_charispd[ii*GT_BYTES+jj]  <= #TCQ 0;
            PPG_gtrx_charissc[ii*GT_BYTES+jj]  <= #TCQ 0;
          end else begin
            PPG_gtrx_charisa[ii*GT_BYTES+jj]   <= #TCQ is_a[jj];
            PPG_gtrx_charisk[ii*GT_BYTES+jj]   <= #TCQ is_k[jj];
            PPG_gtrx_charisr[ii*GT_BYTES+jj]   <= #TCQ is_r[jj];
            PPG_gtrx_charism[ii*GT_BYTES+jj]   <= #TCQ is_m[jj];
            PPG_gtrx_charispd[ii*GT_BYTES+jj]  <= #TCQ is_pd[jj];
            PPG_gtrx_charissc[ii*GT_BYTES+jj]  <= #TCQ is_sc[jj];
          end
        end
      end // end for (jj < GT_BYTES)
    end // end for (ii < LINK_WIDTH)

  //Bypass this extra register if GT_REG is not set.
  end else begin: no_gtreg_gen
    always @(*) begin
      PPG_gtrx_data          = GT_gtrx_data;
      PPG_gtrx_chariskchar   = GT_gtrx_charisk;
      PPG_gtrx_chariscomma   = GT_gtrx_chariscomma;
      PPG_gtrx_invalid       = GT_gtrx_disperr | GT_gtrx_notintable;
      PPG_gtrx_chanisaligned = GT_gtrx_chanisaligned;
      PPG_gtrx_reset_req     = GT_gtrx_reset_req;
      PPG_gtrx_reset_done    = GT_gtrx_reset_done;
    end

    for (ii=0; ii < LINK_WIDTH; ii=ii+1) begin : charisx_gen
      wire [GT_BYTES-1:0] is_k;
      wire [GT_BYTES-1:0] is_r;
      wire [GT_BYTES-1:0] is_m;
      wire [GT_BYTES-1:0] is_pd;
      wire [GT_BYTES-1:0] is_sc;
      wire [GT_BYTES-1:0] is_a;

      for (jj=0; jj < GT_BYTES; jj=jj+1) begin: charisx_gtbytes_gen
        assign is_a[jj] = GT_gtrx_charisk[(ii*GT_BYTES)+jj] & 
                          (GT_gtrx_data[((ii*GT_BYTES*8)+(jj*8))+:8] == A_CHAR);
        assign is_k[jj] = GT_gtrx_charisk[(ii*GT_BYTES)+jj] & 
                          (GT_gtrx_data[((ii*GT_BYTES*8)+(jj*8))+:8] == K_CHAR);
        assign is_r[jj] = GT_gtrx_charisk[(ii*GT_BYTES)+jj] & 
                          (GT_gtrx_data[((ii*GT_BYTES*8)+(jj*8))+:8] == R_CHAR);
        assign is_m[jj] = GT_gtrx_charisk[(ii*GT_BYTES)+jj] & 
                          (GT_gtrx_data[((ii*GT_BYTES*8)+(jj*8))+:8] == M_CHAR);
        assign is_pd[jj] = GT_gtrx_charisk[(ii*GT_BYTES)+jj] & 
                          (GT_gtrx_data[((ii*GT_BYTES*8)+(jj*8))+:8] == PD_CHAR);
        assign is_sc[jj] = GT_gtrx_charisk[(ii*GT_BYTES)+jj] & 
                          (GT_gtrx_data[((ii*GT_BYTES*8)+(jj*8))+:8] == SC_CHAR);

        always @(*) begin
          PPG_gtrx_charisa[ii*jj]   = is_a[jj];
          PPG_gtrx_charisk[ii*jj]   = is_k[jj];
          PPG_gtrx_charisr[ii*jj]   = is_r[jj];
          PPG_gtrx_charism[ii*jj]   = is_r[jj];
          PPG_gtrx_charispd[ii*jj]  = is_pd[jj];
          PPG_gtrx_charissc[ii*jj]  = is_sc[jj];
        end
       
      end // end for (jj < GT_BYTES)
    end // end for (ii < LINK_WIDTH)
  end endgenerate // end if (GT_REG)

endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/phy/oplm/srio_gen2_v4_1_16_oplm_init.v#1 $
//----------------------------------------------------------------------
//
// OPLM_INIT
// Description:
// This module contains all the lane initialization state machines
// needed to bring up the link between the SRIO core and its link partner
// This includes the Lane Sync, Lane Alignment, Mode Detect, and
// initialization state machines.  For further details on the state machines
// functionality see the Physical Layer Specification Section 4.12.
//
// Hierarchy:
// PHY_TOP
//    |___OPLM_TOP
//            |___OPLM_INIT <-- this module
// ---------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_oplm_init
  #(
    parameter TCQ          = 100,
    parameter MODE_XG      = 5,                     // {1, 2, 4}
    parameter LINK_WIDTH   = 1,                     // {1, 2, 4}
    parameter GT_BYTES     = 4,                     // Bytes on the GT Interface
    parameter DATA_WIDTH   = LINK_WIDTH*GT_BYTES*8, // Data width
    parameter CHARIS_WIDTH = LINK_WIDTH*GT_BYTES,   // Charisk bus width
    parameter IDLE1        = 1,                     // {0, 1}
    parameter IDLE2        = 0,                     // {0, 1}
    parameter SIM_TRAIN    = 0)                     // {0: FULL, 1: DIVIDED}  
  (
    // {{{ port declarations ---------------
    // System Signals
    input                             gt_pcs_clk,             //GT Clock
    input                             gt_pcs_rst_q,           //GT Clock Reset
    input                             sim_train_en,           //Enable the SIM_TRAIN parameter

    //User Global
    input                             UG_force_reinit,        //Force link reinit

    //Config Interface
    input   [2:0]                     PC_force_lane,          //Force train down
    input                             PC_port_disable,        //Disable link init.

    //Internal Signals
    output reg                        PPI_mode_1x,            //Mode 1x Selected
    output reg                        PPI_rx_lane_r,          //Mode 1x Selected
    output reg  [LINK_WIDTH-1:0]      PPI_lane_sync,          //Lanes in Sync
    output reg                        PPI_port_initialized,   //Port is Init
    output reg                        PPI_reinit_sm,          //Re-initialize
    output reg                        PPI_idle_select_en,     //Look for the IDLE sequence
    input                             PPR_idle_selected,      //Idle seq is sel
    
    //MGT Interface
    input       [CHARIS_WIDTH-1:0]    PPG_gtrx_charispd,      //Character is /PD/
    input       [CHARIS_WIDTH-1:0]    PPG_gtrx_charissc,      //Character is /SC/
    input       [CHARIS_WIDTH-1:0]    PPG_gtrx_chariscomma,   //Character is Comma
    input       [CHARIS_WIDTH-1:0]    PPG_gtrx_invalid,       //Not in Table
    input       [LINK_WIDTH-1:0]      PPG_gtrx_chanisaligned, //Channel is Aligned
    input       [CHARIS_WIDTH-1:0]    PPG_gtrx_charisa,       //Char is /A/
    input                             PPG_gtrx_reset_req,     //RX Buffer Error
    input       [LINK_WIDTH-1:0]      PPG_gtrx_reset_done,    //RX Buffer Resets Done
    output reg                        PPI_gtrx_reset,         //Reset the RX Buffers
    output reg                        PPI_gtrx_chanbonden,    //En Chanel Bonding
    output reg  [LINK_WIDTH-1:0]      PPI_gttx_inhibit,       //TX inhibit

    //Signals for Debug
    output reg                        PPI_n_lanes_aligned,
    output reg                        PPI_n_lanes_rdy,
    output reg  [3:0]                 PPI_init_state,
    output reg                        PPI_x1_mode_detected
    // }}} end port declarations -----------
  );

  // {{{ Local Parameters ------------------
  // Silence Timeout Values based on the baud rate and SIM parameter
  // For all modes this will timeout at 120 (us)
  localparam SILENCE_TIMEOUT_IMP = (MODE_XG == 1) ? 3750 :
                                   (MODE_XG == 2) ? 7500 :
                                   (MODE_XG == 3) ? 9375 :
                                   (MODE_XG == 5) ? 15000 : 18750;//CR768778 fix

  localparam SILENCE_TIMEOUT_SIM = (MODE_XG == 1) ? 51 :
                                   (MODE_XG == 2) ? 52 :
                                   (MODE_XG == 3) ? 53 :
                                   (MODE_XG == 5) ? 55 : 56;

  // this needs to be a wire since it is gated with sim_train_en. however,
  // sim_train_en will be tied off at the top level
  wire [15:0] SILENCE_TIMEOUT = (sim_train_en) ? SILENCE_TIMEOUT_SIM : 
                                                 SILENCE_TIMEOUT_IMP;

  //Discovery Timeout Values
  //for all modes this will timeout at 28 (ms)
  localparam DISC_TIMEOUT_IMP = (MODE_XG == 1) ? 875000 :
                                (MODE_XG == 2) ? 1750000 :
                                (MODE_XG == 3) ? 2187500 :
                                (MODE_XG == 5) ? 3500000 : 4375000;//CR768778 fix

  localparam DISC_TIMEOUT_SIM_DIV = (MODE_XG == 1) ? 10001 :
                                    (MODE_XG == 2) ? 10002 :
                                    (MODE_XG == 3) ? 10003 :
                                    (MODE_XG == 5) ? 10005 : 10006;

  // this needs to be a wire since it is gated with sim_train_en. however,
  // sim_train_en will be tied off at the top level 
  wire [21:0] DISC_TIMEOUT = (sim_train_en) ? DISC_TIMEOUT_SIM_DIV : 
                                              DISC_TIMEOUT_IMP;                            

  //The Redundancy Lane                               
  localparam R = (LINK_WIDTH == 2) ? 1 : 
                 (LINK_WIDTH == 4) ? 2 : 0;

  //State Machine Count Values
  //V_MAX recomemend counts to 4096, divide this by the number of bytes received per cycle
  localparam V_MAX = 10; //valid char count for implementaton 

  //Similarly for V_MAX_SYNC a recomended value is 255.  For a four byte interface 64 is used.
  //(For here we can just look at the high bit [6])
  localparam V_MAX_SYNC = 6;

  // The dcounter counts the data lanes when using a x2 core. 3 is the recomended initial
  // value
  localparam D_MAX = 3;   

  //For the comma counter the recomemned value is 128 bytes.  Th
  //the k_ctr will count until [K_MAX] is 1.
  localparam K_MAX = 7;

  //Used in the Mode Detect State Machine.
  localparam PD_CHAR = 8'h7C;
  localparam SC_CHAR = 8'h1C;

  //State Machine States
  localparam INIT_SILENT        = 4'd0;
  localparam INIT_SEEK          = 4'd1;
  localparam INIT_SYNC_WAIT     = 4'd2;
  localparam INIT_DISCOVERY     = 4'd3;
  localparam INIT_GTRX_RESET    = 4'd4;
  localparam INIT_NX_MODE       = 4'd5;
  localparam INIT_1X_MODE_LN0   = 4'd6;
  localparam INIT_1X_MODE_LNR   = 4'd7;
  // }}} Local Parameters ------------------

  // {{{ Wire Declarations -----------------
  wire  [GT_BYTES-1:0]        rx_charispd     [LINK_WIDTH-1:0];
  wire  [GT_BYTES-1:0]        rx_charissc     [LINK_WIDTH-1:0];
  wire  [GT_BYTES-1:0]        rx_chariscomma  [LINK_WIDTH-1:0];
  wire  [GT_BYTES-1:0]        rx_invalid      [LINK_WIDTH-1:0];
  reg                         silent_tmr_en;
  reg                         disc_tmr_en;
  reg   [23:0]                tmr;
  reg                         tmr_done;
  reg   [3:0]                 init_next_state;
  reg   [LINK_WIDTH-1:0]      inhibit;
  reg                         idle_select_en;
  reg                         gtrx_reset;
  reg                         rx_lane_r;
  reg                         chanbonden;
  reg                         mode_1x_d;
  reg                         port_init;
  wire                        force_1x;
  wire                        force_lane_r;
  reg   [2:0]                 force_lane_q;
  wire                        force_lane_change;
  // }}} Wire Declarations -----------------
  
  // {{{ if SIMULATION
  //Make State Machine States readable in the waveform
  `ifdef SIMULATION
    reg [20*8-1:0] init_next_state_string = "null";
    reg [20*8-1:0] init_state_string      = "null";

    always @* begin
      case (PPI_init_state)
        INIT_SILENT:      init_state_string = "INIT_SILENT";
        INIT_SEEK:        init_state_string = "INIT_SEEK";
        INIT_SYNC_WAIT:   init_state_string = "INIT_SYNC_WAIT";
        INIT_DISCOVERY:   init_state_string = "INIT_DISCOVERY";
        INIT_GTRX_RESET:  init_state_string = "INIT_GTRX_RESET";
        INIT_NX_MODE:     init_state_string = "INIT_NX_MODE";
        INIT_1X_MODE_LN0: init_state_string = "INIT_1X_MODE_LN0";
        INIT_1X_MODE_LNR: init_state_string = "INIT_1X_MODE_LNR";
        default:          init_state_string = "INVALID";
      endcase
      case (init_next_state)
        INIT_SILENT:      init_next_state_string = "INIT_SILENT";
        INIT_SEEK:        init_next_state_string = "INIT_SEEK";
        INIT_SYNC_WAIT:   init_next_state_string = "INIT_SYNC_WAIT";
        INIT_DISCOVERY:   init_next_state_string = "INIT_DISCOVERY";
        INIT_GTRX_RESET:  init_next_state_string = "INIT_GTRX_RESET";
        INIT_NX_MODE:     init_next_state_string = "INIT_NX_MODE";
        INIT_1X_MODE_LN0: init_next_state_string = "INIT_1X_MODE_LN0";
        INIT_1X_MODE_LNR: init_next_state_string = "INIT_1X_MODE_LNR";
        default:          init_next_state_string = "INVALID";
      endcase
    end
  `endif
  // }}} if SIMULATION
  
  // {{{ MGT Interface ---------------------
  // Split up the MGT signals into a 2-dimentional array for easy access to each
  // lanes values.
  genvar d_ii;
  generate
    //Expand the gtrx_data bus out into a two dimensional array to easily
    //access throughout this module
    for (d_ii = 0; d_ii < LINK_WIDTH; d_ii = d_ii+1) begin: expand_rx_gen
      assign rx_charispd[d_ii]    = PPG_gtrx_charispd[(d_ii*GT_BYTES)+:GT_BYTES];
      assign rx_charissc[d_ii]    = PPG_gtrx_charissc[(d_ii*GT_BYTES)+:GT_BYTES];
      assign rx_chariscomma[d_ii] = PPG_gtrx_chariscomma[(d_ii*GT_BYTES)+:GT_BYTES];
      assign rx_invalid[d_ii]     = PPG_gtrx_invalid[(d_ii*GT_BYTES)+:GT_BYTES];
    end
  endgenerate
  // }}} MGT Interface ---------------------

  // {{{ Lane Synchronization --------------
  // The lane sync state machine counter comma characters, valid code-groups,
  // and invalid code-groups to obtain lane synchronization.  This state
  // machine counter is modeled after Figure 4-4 in the PHY layer
  // specification.
  // There is one lane sync state machine for every lane.

  //These are created outside the scope of the generate in order to assist
  //in coverage in the bind files.  This enables automatic binding and
  //eliminates the need for heirarchical references.
  reg  [7:0]            k_ctr  [LINK_WIDTH-1:0];
  reg  [10:0]           v_ctr  [LINK_WIDTH-1:0];
  reg  [2:0]            i_ctr  [LINK_WIDTH-1:0];
  wire [LINK_WIDTH-1:0] k_ctr_rst;
  wire [LINK_WIDTH-1:0] v_ctr_rst;
  wire [LINK_WIDTH-1:0] i_ctr_rst;
  reg  [LINK_WIDTH-1:0] v_max_pre_sync;

  genvar sync_ii;// lane sync state machine for each lane loop
  //Generate the sync state machine for each lane
  generate 
    for (sync_ii = 0; sync_ii < LINK_WIDTH; sync_ii=sync_ii+1) begin: sync_sm_gen
      wire  lane_synced_aquired;
      reg   first_valid_comma_detect;
      reg   valid_comma_detect;

      // If a valid comma is detected on the same cycle as an invalid we need to
      // detect if it needs to be counted.
      always @* begin
        casex (rx_invalid[sync_ii])
          4'bXXX1: valid_comma_detect = 1'b0;
          4'bXX10: valid_comma_detect = rx_chariscomma[sync_ii][0];
          4'bX100: valid_comma_detect = |rx_chariscomma[sync_ii][1:0];
          4'b1000: valid_comma_detect = |rx_chariscomma[sync_ii][2:0];
          4'b0000: valid_comma_detect = |rx_chariscomma[sync_ii];
          default: valid_comma_detect = 1'bX;
        endcase
      end

      //*COVERAGE*
      // (cp_kcounter_overcount): check that the k gets more commas than needed
      // to reach its max value before it is already maxed
      
      //Comma Counter
      //A comma counter reset should occur if:
      //1. an invalid is detected before sync
      //2. i_ctr reached Imax after sync (after sync is not needed in this
      //expression since the i_ctr only counts after sync).
      assign k_ctr_rst[sync_ii] = (|rx_invalid[sync_ii] & ~PPI_lane_sync[sync_ii]) | 
                                  (i_ctr[sync_ii][2]);

      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          k_ctr[sync_ii] <= #TCQ 0;
        end else begin
          if (!valid_comma_detect && k_ctr_rst[sync_ii]) begin
            k_ctr[sync_ii] <= #TCQ 0;

          // If a reset occurs on the same cycle as a valid comma 
          // Restart with the new comma values
          end else if (k_ctr_rst[sync_ii] && !(k_ctr[sync_ii][K_MAX])) begin
            // But sure the invalid byte is not used to increment with in case
            // it was a "comma"
            casex (rx_invalid[sync_ii])
              //4'bXXX1 will never happen since valid_comma_detect will be
              //0 if rx_invalid is set and the above condition will be entered
              //based on line 247 above
              4'bXX10: begin
                k_ctr[sync_ii] <= #TCQ rx_chariscomma[sync_ii][0];
              end
              4'bX100: begin
                k_ctr[sync_ii] <= #TCQ rx_chariscomma[sync_ii][0] + 
                                       rx_chariscomma[sync_ii][1];
              end
              4'b1000: begin
                k_ctr[sync_ii] <= #TCQ rx_chariscomma[sync_ii][0] + 
                                       rx_chariscomma[sync_ii][1] + 
                                       rx_chariscomma[sync_ii][2];
              end
              default: k_ctr[sync_ii] <= #TCQ {LINK_WIDTH{1'bX}};
            endcase

          // else Increment                       
          end else if (!(k_ctr[sync_ii][K_MAX])) begin
            k_ctr[sync_ii] <= #TCQ k_ctr[sync_ii] + rx_chariscomma[sync_ii][0] + 
                                                    rx_chariscomma[sync_ii][1] +
                                                    rx_chariscomma[sync_ii][2] +
                                                    rx_chariscomma[sync_ii][3];
          end
        end
      end

      //*COVERAGE*
      //(cp_comma_counts): See all possible counters of comma characters arrive for the 
      // K counter before it is maxed
 
      //Valid Code-groups Counter
      //A valid rest should occur if:
      //1. An invalid byte is detected
      //2. i_ctr reaches i_max (4)
      //4. lane sync is reached and we can now start after sync counter
      //5. The first valid comma is not yet found.
      assign v_ctr_rst[sync_ii] = |rx_invalid[sync_ii] | i_ctr[sync_ii][2] | 
                                  lane_synced_aquired  | !first_valid_comma_detect;



      // The valid codegroups counter should start counting after the first
      // valid comma is detected
      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          first_valid_comma_detect <= #TCQ 0;
        end else begin
          if (!valid_comma_detect && k_ctr_rst[sync_ii]) begin
            first_valid_comma_detect <= #TCQ 0;
          end else if (|rx_chariscomma[sync_ii]) begin
            first_valid_comma_detect <= #TCQ 1;
          end
        end
      end

      // Count the valid codegroups when not in a counter reset state
      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          v_max_pre_sync[sync_ii] <= #TCQ 0;
        end else begin
          if (v_ctr_rst[sync_ii]) begin
            v_max_pre_sync[sync_ii] <= #TCQ 0;
          end else if ((v_ctr[sync_ii][V_MAX]) && !PPI_lane_sync[sync_ii]) begin
            v_max_pre_sync[sync_ii] <= #TCQ 1;
          end
        end
      end

      //*COVERAGE*
      //(cp_vcounter_reset_pre_sync): See the v counter reset before lane sync

      //*COVERAGE*
      //(cp_vcounter_reset_post_sync): See the v counter reset after lane sync

      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          v_ctr[sync_ii] <= #TCQ 0;
        end else begin
          if (v_ctr_rst[sync_ii]) begin
            v_ctr[sync_ii] <= #TCQ 0;

          end else begin
            //Increment the counter for every valid four bytes detected. 
            //This counter is free running unless a reset condition occurs.
            v_ctr[sync_ii] <= #TCQ v_ctr[sync_ii] + 1'b1;
          end
        end
      end

      //*COVERAGE*
      //(cp_vcounter_rollsover): See the v counter roll over

      //*COVERPOINT*
      // (cp_lane_sync): All combinations of lane synchronization are hit to varify 
      // that lanes come up in various orders and the redundancy lane is used.
  
      assign lane_synced_aquired = v_max_pre_sync[sync_ii] && k_ctr[sync_ii][K_MAX];

      //Drive the lane sync signal
      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          PPI_lane_sync[sync_ii] <= #TCQ 0;
        end else begin
          //The lane is in sync
          if (lane_synced_aquired) begin
            PPI_lane_sync[sync_ii] <= #TCQ 1'b1;

          //When the invalid counter reaches it max the lane is no longer in
          //sync
          end else if (i_ctr[sync_ii][2]) begin
            PPI_lane_sync[sync_ii] <= #TCQ 1'b0;
          end
        end
      end

      //Invalid Code-groups Counter
      //This counter should hold a value of 0 as long as the lane is not in
      //sync.
      assign i_ctr_rst[sync_ii] = (!PPI_lane_sync[sync_ii]) | (i_ctr[sync_ii][2]);

      //*ASSERTION*
      //(ap_icounter_rollunder): i_ctr (invalid code-groups) decrements to past 0

      //*COVERPOINT*
      //(cp_icounter_max): The Invalid code groups counter finds its max value of 
      // 4 invalid groups
      
      //*ASSERTION*
      //(ap_icounter_rollover): The i_ctr must not roll over the max value of 7

      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          i_ctr[sync_ii] <= #TCQ 0;
        end else begin
          if (i_ctr_rst[sync_ii]) begin
            i_ctr[sync_ii] <= #TCQ 0;

          //Increment the counter for any invalid byte detected
          end else if (|rx_invalid[sync_ii] && !i_ctr[sync_ii][2]) begin
            i_ctr[sync_ii] <= #TCQ i_ctr[sync_ii] + rx_invalid[sync_ii][0] + rx_invalid[sync_ii][1] +
                                                    rx_invalid[sync_ii][2] + rx_invalid[sync_ii][3];

          //After sync is obtained, decrement the invalid count if there was
          //v_max number of valid bytes detected since the last invalid byte
          end else if (PPI_lane_sync[sync_ii] && (i_ctr[sync_ii] > 0) && (v_ctr[sync_ii][V_MAX_SYNC])) begin
            i_ctr[sync_ii] <= #TCQ i_ctr[sync_ii] - 1'b1;
          end
        end
      end
    end //end for (sync_ii < LINK_WIDTH)
  endgenerate
  // }}} Lane Synchronization --------------

  // {{{ Lane Alignment --------------------
  // The lane alignment state machine monitors the alignment of data through
  // the MGTs.  This state machine is modeled after Figure 4-15 of the PHY
  // layer specification.  This is only required for multii-lane
  // configurations.

  //These are created outside the scope of the generate in order to assist
  //in coverage in the bind files.  This enables automatic binding and
  //eliminates the need for heirarchical references.
  //The max value of the a and m counter are 4 as indicated in the PHY
  //layer spec section 4.12.4.3
  reg   [2:0]           a_ctr;
  reg   [2:0]           m_ctr;
  wire                  a_ctr_rst;
  wire                  m_ctr_rst;
  wire  [GT_BYTES-1:0]  misaligned_column;
  wire  [GT_BYTES-1:0]  a_column;
  wire  [GT_BYTES-1:0]  a_detect;
  genvar                a_ii;   // a char expand
  genvar                acb_ii; // a columns bytes
  genvar                ma_ii;  // miasligned a count 

  //Generate the lane alignment state machine when the link width is 
  //greater than 1. Otherwise, tie of the PPI_n_lanes_aligned output
  //to not interfer with the initialization state machine.
  generate
    if (LINK_WIDTH > 1) begin: lane_align_sm_gen

      wire [GT_BYTES-1:0] charisa  [LINK_WIDTH-1:0];
      
      for (a_ii=0; a_ii < LINK_WIDTH; a_ii=a_ii+1) begin: a_expand_gen
        assign charisa[a_ii] = PPG_gtrx_charisa[a_ii*GT_BYTES+:GT_BYTES];
      end

      if (LINK_WIDTH == 2) begin: x2_a_gen
        for (acb_ii=0; acb_ii < GT_BYTES; acb_ii=acb_ii+1) begin: a_col_det_gen
          assign a_column[acb_ii] = charisa[0][acb_ii] & charisa[1][acb_ii];
          assign a_detect[acb_ii] = charisa[0][acb_ii] | charisa[1][acb_ii];
        end

      end else if (LINK_WIDTH == 4) begin: x4_a_gen
        for (acb_ii=0; acb_ii < GT_BYTES; acb_ii=acb_ii+1) begin: a_col_det_gen
          assign a_column[acb_ii] = charisa[0][acb_ii] & charisa[1][acb_ii] & 
                                    charisa[2][acb_ii] & charisa[3][acb_ii];
          assign a_detect[acb_ii] = charisa[0][acb_ii] | charisa[1][acb_ii] | 
                                    charisa[2][acb_ii] | charisa[3][acb_ii];
        end
      end

      //"A" Character Counter
      //Counts the number of columns of "A"s.
      //A reset occurs if:
      //1. all the lanes are not in sync
      //2. the m_ctr has started counting
      //3. the a_ctr reaches its max and n_lanes_aligned is going to assert
      //4. a misalignment is detected
      assign a_ctr_rst = ~(&PPI_lane_sync) || (PPI_n_lanes_aligned && (m_ctr == 0)) || 
                          a_ctr[2]         || (|misaligned_column);

      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          a_ctr <= #TCQ 0;
        end else begin
          if (a_ctr_rst) begin
            a_ctr <= #TCQ 0;

          // Increment for every a column detected
          end else begin
            a_ctr <= #TCQ a_ctr + a_column[0] + a_column[1] + a_column[2] + a_column[3];
          end
        end
      end

      //*ASSERTION*
      //(ap_acounter_underflow): Alignment counter does not underflow

      //*ASSERTION*
      //(ap_acounter_rollover): The a_ctr must not roll over the max value of 7

      //*COVERAGE*
      //(cp_a_column): Cover all interesting values of a_column

      //*COVERAGE*
      //(cp_a_detect): Cover all interesting values of a_detect when there is
      //not a column of A's

      //*COVERPOINT*
      //(cp_acounter_max): The Alignment counter reaches its max value

      //*COVERPOINT*
      //(cp_align_err_before_aligned): before alignment is obtain, an alignment 
      // error is seen

      //*COVERPOINT*
      //(cp_align_err_after_aligned): and alignment error is seen after alignment
      // is obtained

      //Drive PPI_n_lanes_aligned
      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          PPI_n_lanes_aligned <= #TCQ 1'b0;
        end else begin
          if (~(&PPI_lane_sync) || m_ctr[2])
            PPI_n_lanes_aligned <= #TCQ 1'b0;
          else if (a_ctr[2])
            PPI_n_lanes_aligned <= #TCQ 1'b1;
        end
      end

      //Misalignment Counter
      //Counts the number of times it sees a misaligned colum after
      //PPI_n_lanes_aligned is asserted.
      //If the max number of |A|'s are seen before the m counter maxes,
      //reset the count.
      assign m_ctr_rst = ~(PPI_n_lanes_aligned) || a_ctr[2];

      //A column is missagligned if an A is seen but it is not
      //across all the lanes.
      for (ma_ii=0; ma_ii < GT_BYTES; ma_ii=ma_ii+1) begin: misaligned_a_gen
        assign misaligned_column[ma_ii] = a_detect[ma_ii] && !a_column[ma_ii];
      end

      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          m_ctr <= #TCQ 0;
        end else begin
          if (m_ctr_rst) begin
            m_ctr <= #TCQ 0;
          end else begin
            m_ctr <= #TCQ m_ctr + misaligned_column[0] + misaligned_column[1]  + 
                                  misaligned_column[2] + misaligned_column[3];
          end
        end
      end
      //*ASSERTION*
      //(ap_mcounter_rollover): The m_ctr must not roll over the max value of 7

      //*COVERPOINT*
      //(cp_mcounter_max): The misalignement counter reaches its max value
      // after PPI_n_lanes_aligned was asserted
      
      //*COVERAGE*
      //(cp_misaligned_column): cover a misaligned column is seen in each byte
      // location
    end //end if (LINK_WIDTH > 1)
    else begin: lane_align_1x_gen
      // For 1x cores, the PPI_n_lanes_aligned signal is always asserted
      // for use in the initialization state machine
      always @(posedge gt_pcs_clk) begin
        PPI_n_lanes_aligned <= #TCQ 1'b0;
      end
    end
  endgenerate
  // }}} Lane Alignment --------------------

  // {{{ Mode Detect (2x Only) -------------
  //These are created outside the scope of the generate in order to assist
  //in coverage in the bind files.  This enables automatic binding and
  //eliminates the need for heirarchical references.
  reg [1:0]   d_ctr;
  wire        x1_mode_delimit;
  wire        x2_mode_delimit;
  wire        d_ctr_rst;

  //Generate the mode detection state machine only when the link width is 2x.
  //Otherwise tie off the PPI_x1_mode_detected signal output to not interfer with 
  //the initialization state machine.
  genvar md_ii; //mode delimit
  generate 
    if (LINK_WIDTH == 2) begin: mode_detect_sm_gen
      // The mode detect state machine determines if a 2x cores is in 1x mode
      // or 2x mode. This models the state machine in Figure 4-16 of the PHY
      // layer specification.
      wire                pdsc_laner_byte0;
      wire                pdsc_lane0_byte1;
      wire                pdsc_laner_byte1;
      reg                 n_lanes_aligned_q;
      wire [GT_BYTES-1:0] x1_mode_delimit_d;
      wire [GT_BYTES-1:0] x2_mode_delimit_d;

      //Monitor for a change in PPI_n_lanes_aligned
      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          n_lanes_aligned_q <= #TCQ 0; 
        end else begin
          n_lanes_aligned_q <= #TCQ PPI_n_lanes_aligned;
        end
      end

      //*COVERPOINT*
      //(cp_x1_mode_delimit): A x2 is recognized as in x1 mode
     
      //*COVERPOINT*
      //(cp_x2_mode_delimit): A x2 is recognized as in x2 mode

      for (md_ii=0; md_ii < GT_BYTES; md_ii=md_ii+1) begin: mode_delimit_gen
        /// Receiving in 1x mode if a PD/SC is on both lanes on the same byte
        assign x1_mode_delimit_d[md_ii] = (rx_charispd[R][md_ii] || rx_charissc[R][md_ii]) && 
                                          (rx_charispd[0][md_ii] || rx_charissc[0][md_ii]);

        // Receiving in 2x mode if a PD/SC is only seen on one lane on a given byte
        assign x2_mode_delimit_d[md_ii] = (rx_charispd[0][md_ii] ^ rx_charissc[R][md_ii]) ||
                                          (rx_charispd[0][md_ii] ^ rx_charissc[R][md_ii]);
      end
      assign x1_mode_delimit = |x1_mode_delimit_d;
      assign x2_mode_delimit = |x2_mode_delimit_d;

      //The D counter is an up/down counter to monitor the state of the lanes
      //for a 2x core.  
      //A reset occurs if there is a change in the lanes alignment
      assign d_ctr_rst = (n_lanes_aligned_q != PPI_n_lanes_aligned) | ~(PPI_n_lanes_aligned);
                       
      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          d_ctr <= #TCQ D_MAX;
        end else begin
          if (d_ctr_rst) begin
            d_ctr <= #TCQ D_MAX;

          //only decrement if we are not already 0
          end else if (x1_mode_delimit && (|d_ctr)) begin
            d_ctr <= #TCQ d_ctr - 1;

          //Only increment if we are not at the max value
          end else if (x2_mode_delimit && !(&d_ctr)) begin
            d_ctr <= #TCQ d_ctr + 1;
          end
        end
      end
      
      //*ASSERTION*
      //(ap_dcounter_underflow): Check that the d_ctr does not underflow

      //*ASSERTION*
      //(ap_dcounter_overflow): Check that the d_ctr does not overflow

      // Assert 1x mode once the d_ctr gets to 0
      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          PPI_x1_mode_detected <= #TCQ 1'b0;
        end else begin
          if (d_ctr_rst) begin
            PPI_x1_mode_detected <= #TCQ 1'b0;

          end else if (d_ctr == 0) begin 
            PPI_x1_mode_detected <= #TCQ 1'b1;
          end
        end
      end

      //*COVERAGE*
      //(cp_dcounter_reached_zero):  The d counter reaches 0 and a x2 is now
      // in x1 mode.

    end //end if (LINK_WIDTH == 2)
    else begin: no_mode_det_sm_gen
      //Tire the 1x mode detected signal low for other link widths.
      //1x mode will be detemined by the initialization state machine.
      always @(posedge gt_pcs_clk) begin
        PPI_x1_mode_detected <= #TCQ 1'b0;
      end
    end
  endgenerate
  // }}} Mode Detect (2x Only) -------------

  // {{{ Initialization --------------------
  //Timer to calculate how long to stay in the silent and discovery states
  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      tmr <= #TCQ 0;
    end else begin
      //If no timer is enabled, or a state machine reinit occurs, reset
      if ((!silent_tmr_en && !disc_tmr_en) || PPI_reinit_sm) begin
        tmr <= #TCQ 0;
      end else begin
        //Only count until the max value is reached.
        if (!(tmr_done))
          tmr <= #TCQ tmr + 1'b1;
      end
    end
  end

  //Register if the timer has reaches it max count value
  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      tmr_done <= #TCQ 0; 
    end else begin
      if (PPI_reinit_sm) begin
        tmr_done <= #TCQ 0;
      end else begin
        tmr_done <= #TCQ (silent_tmr_en & (tmr >= SILENCE_TIMEOUT)) |
                         (disc_tmr_en   & (tmr >= DISC_TIMEOUT));
      end
    end 
  end

  //all the lanes are ready if they are all in sync and aligned
  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      PPI_n_lanes_rdy <= #TCQ 0;
    end else begin
      PPI_n_lanes_rdy <= #TCQ &PPI_lane_sync & PPI_n_lanes_aligned;
    end
  end

  //*COVERPOINT*
  //(cp_Nx_not_rdy_no_sync): In xN mode with the port initialized, PPI_n_lanes_rdy 
  // is deasserted with sync on no lanes.
  
  //*COVERPOINT*
  //(cp_Nx_not_rdy_sync): In xN mode with the port initialized, PPI_n_lanes_rdy 
  // is deasserted with sync on a lane.

  //Register the force_lane signal to reinit the state machine if it updates
  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      force_lane_q <= #TCQ 0;
    end else begin
      force_lane_q <= #TCQ PC_force_lane;
    end
  end

  assign force_lane_change = force_lane_q != PC_force_lane;

  //Force x1 conditions
  assign force_1x     = (PC_force_lane == 3'b010) || (PC_force_lane == 3'b011); 
  assign force_lane_r = (PC_force_lane == 3'b011);
    
  //Create this local parameter only used in this state machine to by pass
  //warnings generated by vsim. This signal is only used when LINK_WIDTH == 4
  //to disable lanes 1 and 3 when the core is trained to 1x.
  localparam LANE1 = (LINK_WIDTH == 4) ? 1 : 0;
  localparam LANE3 = (LINK_WIDTH == 4) ? 3 : 0;

  //Wires used to simplify the condition for INIT_DISCOVERY -> INIT_1X_MODE_LN0
  wire force_lane_r_failed = force_1x && force_lane_r && tmr_done && !PPI_lane_sync[R];
  wire force_lane0         = force_1x && !force_lane_r;
  wire lanes_not_rdy0      = !force_lane_r && tmr_done && !PPI_n_lanes_rdy;
  wire x2_resolved_as_x1   = PPI_n_lanes_rdy && PPI_x1_mode_detected;

  //Wires used to simplify the condition for INIT_DISCOVERY -> INIT_1X_MODE_LNR
  wire forced_lane_r      = force_1x && force_lane_r;
  wire force_lane0_failed = force_1x && !force_lane_r && tmr_done && !PPI_lane_sync[0];
  wire lanes_not_rdy_r    = tmr_done && !PPI_lane_sync[0] && !force_1x && !PPI_n_lanes_rdy;

  always @(*) begin
    //Set Initial defaults
    silent_tmr_en     = 0;
    disc_tmr_en       = 0;
    port_init         = 0;
    rx_lane_r         = 0; 
    gtrx_reset        = 0;
    chanbonden        = 0;
    mode_1x_d         = (LINK_WIDTH == 1);
    idle_select_en    = 0;

    case (PPI_init_state)
      //Disable all output drivers forcing the link partner to reinitialize
      //Remain in the silent state for +/- 40 us.  
      INIT_SILENT: begin
        silent_tmr_en  = 1;
        inhibit        = {LINK_WIDTH{1'b1}};

        if (tmr_done) begin
          init_next_state = INIT_SEEK;
        end else begin
          init_next_state = INIT_SILENT;
        end
      end

      //Turn on lanes 0 and R of the MGTs. Once sync is obtained on at least
      //one lane and the IDLE sequence is known, go to the sync wait state.
      //If its a 1x core and sync is obtained, go directly to the 1x mode
      //state.
      INIT_SEEK: begin
        //Inhibit all the GTs except lanes 0 and R
        inhibit        = {LINK_WIDTH{1'b1}};
        inhibit[0]     = 1'b0;
        inhibit[R]     = 1'b0; //R is 0 w/LINK_WIDTH==1 so no harm in turn it on all the time
        idle_select_en = 1; 

        // On RX buffer errors from the MGTS reset the buffers.
        // Note: This does not wait for reset done, reset done is a pcs reset
        // indicator, there is no indication of completion for a buffer reset
        if (PPG_gtrx_reset_req) begin
          gtrx_reset      = 1'b1;
          init_next_state = INIT_SEEK;

          //*COVERPOINT*
          //(cp_resetreq_from_seek): A RX buf error occurs in the seek state
        end else if ((PPI_lane_sync[0] || PPI_lane_sync[R]) && 
                     PPR_idle_selected && (LINK_WIDTH != 1) && !force_1x) begin
          init_next_state = INIT_SYNC_WAIT;
        end else if ((PPI_lane_sync[0] || PPI_lane_sync[R]) && 
                     PPR_idle_selected && (LINK_WIDTH != 1) && force_1x) begin
          init_next_state = INIT_DISCOVERY;
        end else if (PPI_lane_sync[0] && PPR_idle_selected && (LINK_WIDTH == 1)) begin
          init_next_state = INIT_1X_MODE_LN0;
        end else begin
          init_next_state = INIT_SEEK;
        end
      end

      //The Sync wait state waits until all N lanes are in sync and then
      //resets all the RX buffers in the MGTs.  This is required by the GTs in
      //order for then to align/chanel bond properly. This is "a part of the
      //discovery state" and so the discovery timer must start the timer here.
      INIT_SYNC_WAIT: begin
        disc_tmr_en = 1'b1;

        //Enable all the GTs, any that resolve to unused will be turned off
        //when the port initializes
        if (!force_1x) begin
          inhibit = {LINK_WIDTH{1'b0}};
        end else begin
          inhibit = PPI_gttx_inhibit;
        end

        // On RX buffer errors from the MGTS reset the buffers.
        // Note: This does not wait for reset done, reset done is a pcs reset
        // indicator, there is no indication of completion for a buffer reset
        if (PPG_gtrx_reset_req) begin
          gtrx_reset      = 1'b1;
          init_next_state = INIT_SYNC_WAIT;

          //*COVERPOINT*
          //(cp_resetreq_from_sync_wait): A RX buf error occurs in the sync
          // wait state

        end else if (&PPI_lane_sync) begin
          gtrx_reset      = 1'b1;
          init_next_state = INIT_GTRX_RESET;
            
          //*ASSERTION*
          //(ap_bufrst_first_sync): The first lane sync across N lanes issues a buffer reset
          
        end else if (tmr_done) begin
          init_next_state = INIT_DISCOVERY;

          //*COVERPOINT*
          //(cp_to_sync): The discovery timer times out in the init_sync_state
        end else begin
          init_next_state = INIT_SYNC_WAIT;
        end
      end

      //Entering this state mean the rx buffers was reset in the MGTs and we
      //now need to wait till sync is obtained again.  This state is "part of
      //discovery" and must enable the discovery timer.
      INIT_GTRX_RESET: begin
        //*COVERPOINT*
        //(cp_resetreq_from_disc): the INIT_GTRX_RESET state is entered from INIT_DISCOVERY

        disc_tmr_en = 1'b1;

        //Enable all the GTs, any that resolve to unused will be turned off
        //when the port initializes
        if (!force_1x) begin
          inhibit = {LINK_WIDTH{1'b0}};
        end else begin
          inhibit = PPI_gttx_inhibit;
        end
        
        // On RX buffer errors from the MGTS reset the buffers.
        // Note: This does not wait for reset done, reset done is a pcs reset
        // indicator, there is no indication of completion for a buffer reset
        if (PPG_gtrx_reset_req) begin
          gtrx_reset      = 1'b1;
          init_next_state = INIT_GTRX_RESET;

          //*COVERPOINT*
          //(cp_resetreq_from_gtrx_reset): A RX buf error occurs in the
          //gtrx_reset state 
        
          // Do not include coverage for tmr_done asserting in this state since
        // this will never happen in hardware. If there is sync then there
        // should always be a reset_done assertion to follow. If reset done
        // never asserts a hard reset will need to be used to fix the GTs.

        // Note: This waits for reset_done since that is what we validated
        // with and it seemed risky to change it. This in theory should not
        // need to wait for reset done, just sync before going into discovery
        end else if ((PPI_lane_sync[0] && PPG_gtrx_reset_done[0]) || 
                     (PPI_lane_sync[R] && PPG_gtrx_reset_done[R]) || tmr_done) begin
          init_next_state = INIT_DISCOVERY;
            
          //*COVERPOINT*
          //(cp_sync_in_bufrst): Lane sync is seen from the GTRX_RESET state

        end else begin 
          init_next_state = INIT_GTRX_RESET;
        end
      end

      //Stay in the discovery state for 28 +/- 4 msec as indicated by the PHY
      //spec (4.12.4.1.3).  In this state chanel bonding of the MGTs should be
      //enabled when all N lanes are in sync. 
      INIT_DISCOVERY: begin
        disc_tmr_en  = 1'b1;
        chanbonden   = &PPI_lane_sync;

        //Enable all the GTs, any that resolve to unused will be turned off
        //when the port initializes
        if (!force_1x) begin
          inhibit = {LINK_WIDTH{1'b0}};
        end else begin
          inhibit = PPI_gttx_inhibit;
        end

        // On RX buffer errors from the MGTS reset the buffers.
        // Note: This goes into gtrx_reset state and waits for reset_done since 
        // that is what we validated with and it seemed risky to change it. 
        // This in theory should not need to wait for reset done, just assert
        // reset and remain in discovery
        if (PPG_gtrx_reset_req) begin
          gtrx_reset      = 1'b1;
          init_next_state = INIT_GTRX_RESET;

          //*COVERPOINT*
          //(cp_resetreq_from_disc): gtrx_reset_req asserts in the discovery state
          //*ASSERTION*
          //(ap_err_bufrst): An GT RX Buffer Error issues a GT RX Buffer Reset

        //If there is no sync of either lane for 1x mode and the discover
        //timer is done, start back in the silent state.
        end else if ((!PPI_lane_sync[0] && !PPI_lane_sync[R]) && tmr_done) begin
          init_next_state = INIT_SILENT;

          //*COVERPOINT*
          //(cp_to_disc): The discovery timer times out in the discovery state 

        //Initialize to 1x on lane 0 if:
        //1. Forcing 1x to lane 0 is requested and sync was on lane 0
        //2. Force to lane R was request but not achieved, and lane 0 was in
        //   sync when the timer was done
        //3. Not all lanes were rdy for Nx mode when the timer was done, but
        //   lane 0 was in sync.
        //4. for 2x cores, all lanes were rdy and we detected 1x mode. from
        //   monitoring lane 0 and R.
        end else if (PPI_lane_sync[0] && 
                    (force_lane0 || force_lane_r_failed || lanes_not_rdy0 || x2_resolved_as_x1)) begin
          init_next_state = INIT_1X_MODE_LN0;
        
        //Initialize to 1x on lane R if:
        //1. We are forcing lane R init and sync is valid on that lane
        //2. All lanes did not sync by the end of the discovery timer but lane
        //   R has sync and lane 0 does not
        //3. We wanted to force 1x mode to lane 0, but lane 0 did not sync and
        //   lane R did, so just use lane R.
        end else if (PPI_lane_sync[R] && (forced_lane_r || force_lane0_failed || lanes_not_rdy_r)) begin
          init_next_state = INIT_1X_MODE_LNR;  

        //If All lanes are up and we are not forcing a 1x mode the port should
        //initialize.
        end else if (!force_1x && PPI_n_lanes_rdy) begin
          init_next_state = INIT_NX_MODE;

        end else begin
          init_next_state = INIT_DISCOVERY;
        end
      end

      //The port is init to Nx mode
      INIT_NX_MODE: begin
        port_init = 1'b1;

        //Enable all the GTs, any that resolve to unused will be turned off
        //when the port initializes
        inhibit = {LINK_WIDTH{1'b0}};

        if ((!PPI_n_lanes_rdy && (PPI_lane_sync[0] || PPI_lane_sync[R])) || 
            (PPI_n_lanes_rdy && PPI_x1_mode_detected))
          init_next_state = INIT_DISCOVERY;
        else if (!PPI_n_lanes_rdy && !PPI_lane_sync[0] && !PPI_lane_sync[R])
          init_next_state = INIT_SILENT;
        else
          init_next_state = INIT_NX_MODE;
      end

      //The port is init to 1x mode with lane 0 as the primary lane.
      INIT_1X_MODE_LN0: begin
        port_init = 1'b1;
        mode_1x_d = 1'b1;
        inhibit   = {LINK_WIDTH{1'b0}};

        //Disable the MGTs not in use.
        if (LINK_WIDTH == 4) begin
          inhibit[LANE1] = 1'b1;
          inhibit[LANE3] = 1'b1;
        end

        if (!PPI_lane_sync[0])
          init_next_state = INIT_SILENT;
        else
          init_next_state = INIT_1X_MODE_LN0;
      end

      //The port is init to 1x mode with lane R as the primary lane.
      INIT_1X_MODE_LNR: begin
        port_init  = 1'b1;
        mode_1x_d  = 1'b1;
        rx_lane_r  = 1'b1;
        inhibit    = {LINK_WIDTH{1'b0}};

        //Disable the MGTs not in use.
        if (LINK_WIDTH == 4) begin
          inhibit[LANE1] = 1'b1;
          inhibit[LANE3] = 1'b1;
        end 

        if (!PPI_lane_sync[R])
          init_next_state = INIT_SILENT;
        else
          init_next_state = INIT_1X_MODE_LNR;
      end

      default: begin
        silent_tmr_en   = 1'bX;
        disc_tmr_en     = 1'bX;
        port_init       = 1'bX;
        mode_1x_d       = 1'bX;
        rx_lane_r       = 1'bX; 
        gtrx_reset      = 1'bX;
        chanbonden      = 1'bX;
        inhibit         = {LINK_WIDTH{1'b1}};
        idle_select_en  = 1'bX;
        init_next_state = INIT_SILENT;
      end
    endcase
  end

  //Assign outputs based on the init state machine logic
  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      PPI_port_initialized <= #TCQ 0;
    end else begin
      PPI_port_initialized <= #TCQ port_init;
    end
  end

  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      PPI_mode_1x <= #TCQ (LINK_WIDTH == 1);
    end else begin
      PPI_mode_1x <= #TCQ mode_1x_d;
    end
  end

  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      PPI_rx_lane_r <= #TCQ 0;
    end else begin
      PPI_rx_lane_r <= #TCQ rx_lane_r;
    end
  end

  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      PPI_gtrx_reset <= #TCQ 0;
    end else begin
      PPI_gtrx_reset <= #TCQ gtrx_reset;
    end
  end

  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      PPI_gttx_inhibit <= #TCQ -1; //Assign to all 1's
    end else begin
      PPI_gttx_inhibit <= #TCQ inhibit;
    end
  end

  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      PPI_idle_select_en <= #TCQ 0;
    end else begin
      if (PPI_reinit_sm) begin
        PPI_idle_select_en <= #TCQ 0;
      end else begin
        PPI_idle_select_en <= #TCQ idle_select_en;
      end
    end
  end

  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      PPI_gtrx_chanbonden <= #TCQ 0;
    end else begin
      PPI_gtrx_chanbonden <= #TCQ chanbonden;
    end
  end

  //Force a reinitialization of the init state machine by going to SILENT if:
  //1. a force_reinit is issued
  //2. force_lane is written to in the phy cfg regs
  //3. the port is disabled (in which case do not leave the silent state)

  // synchronize the user signal first
  reg [1:0] ug_force_reinit_sync;
  reg       ug_force_reinit_sync_q;
  always @(posedge gt_pcs_clk or posedge UG_force_reinit) begin
    if (UG_force_reinit) begin
      ug_force_reinit_sync <= #TCQ 2'b11;
    end else begin
      ug_force_reinit_sync <= #TCQ {ug_force_reinit_sync[0], 1'b0};
    end
  end

  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      ug_force_reinit_sync_q <= #TCQ 0;
      PPI_reinit_sm          <= #TCQ 0;
    end else begin
      ug_force_reinit_sync_q <= #TCQ |ug_force_reinit_sync;
      PPI_reinit_sm          <= #TCQ ug_force_reinit_sync_q || PC_port_disable || force_lane_change;
    end
  end
  //*COVERPOINT*
  //(cp_reinit_before_init): reinit is forced before PPI_port_initialized
  //(cp_reinit_after_init): reinit is forced after PPI_port_initialized

  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      PPI_init_state <= #TCQ INIT_SILENT;
    end else begin
      if (PPI_reinit_sm)
        PPI_init_state <= #TCQ INIT_SILENT;
      else
        PPI_init_state <= #TCQ init_next_state;
    end
  end
  // }}} Initialization --------------------

 endmodule
// {{{ DISCLAIMER OF LIABILITY
//----------------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/phy/oplm/srio_gen2_v4_1_16_oplm_tx.v#3 $
//----------------------------------------------------------------------
//
// OPLM_TX
// Description:
// This module contains the logic for the TX path of the OPLM.  The TX
// path is responsible for the following:
// 1. Striping any valid data only before transmition
// 2. Generating the appropriate IDLE Sequence
// 3. Generating the Synchronization Sequence if in IDLE2 mode
// 4. Scrambling data prior to transmision 
// 5. Providing this data the GTs to transmit
//
// Hierarchy:
// PHY_TOP
//    |___OPLM_TOP
//            |___OPLM_TX <-- this module
//                    |__EVAL_GT_PCS_CLK
// ---------------------------------------------------------------------
`timescale 1ps/1ps

// ------------------------------------------------
// below attribute is added to supress the synthesis warnings in vivado tool 8:3332
(* DowngradeIPIdentifiedWarnings="yes" *)
// ------------------------------------------------

module srio_gen2_v4_1_16_oplm_tx
  #(
    parameter TCQ           = 100,
    parameter LINK_WIDTH    = 1,                     // {1, 2, 4}
    parameter GT_BYTES      = 4,                     // GT Interface Bytes
    parameter DATA_WIDTH    = LINK_WIDTH*GT_BYTES*8, // Data width
    parameter CHARIS_WIDTH  = LINK_WIDTH*GT_BYTES,   // Charisk bus width
    parameter IDLE1         = 1,                     // {0, 1}
    parameter IDLE2         = 0,                     // {0, 1}
    parameter MODE_XG       = 5,                     // {1, 2, 3, 5, 6}
    parameter SCRAM         = 0,                     // {0, 1}  
    parameter EVAL          = 1)                     // Includes the evaluation timer
  (
    // {{{ port declarations ----------------
    // System Signals
    input                         gt_pcs_clk,          //GT Clock
    input                         gt_pcs_rst_q,        //GT Clock Reset
    input                         phy_clk,              //Phy Clock 
    input                         phy_rst_q,            //Phy Reset 

    // OPLM Synchronization Interface
    input       [63:0]            PT_tx_data,           //Transmit data
    input       [7:0]             PT_tx_charisk,        //Character is K
    input       [1:0]             PT_tx_valid,          //Valid
    input                         PT_tx_early_lreq,     //Clk Comp Granted
    input                         PT_ccomp_grant,       //Clk Comp Granted
    input                         PT_send_lreq,         //Link Request
    output reg                    PPT_lreq_sent,        //Link Request Done
    output reg                    PPT_ccomp_req,        //Clk Comp Request

    // MGT TX Interface
    output reg  [DATA_WIDTH-1:0]  PPT_gttx_data,         //Transmit Data 
    output reg  [CHARIS_WIDTH-1:0]PPT_gttx_charisk,      //Character is K
   
    // PHY Equalization Interface
    input   [LINK_WIDTH-1:0]      PE_gttx_cmd,            // Command to send in the CSF
    input   [LINK_WIDTH*2-1:0]    PE_gttx_tap_m1_cmd,     // Tap -1 Command
    input   [LINK_WIDTH*2-1:0]    PE_gttx_tap_p1_cmd,     // Tap +1 Command
    input   [LINK_WIDTH-1:0]      PE_gttx_reset_emphasis, // Cmd Reset Emphasis
    input   [LINK_WIDTH-1:0]      PE_gttx_preset_emphasis,// Cmd Preset Emphasis
    input   [LINK_WIDTH*2-1:0]    PE_gttx_tap_m1_status,  // Current Tap -1 Status
    input   [LINK_WIDTH*2-1:0]    PE_gttx_tap_p1_status,  // Current Tap +1 Status
    input   [LINK_WIDTH-1:0]      PE_gttx_ack,            // Recieved cmd was ACK'd
    input   [LINK_WIDTH-1:0]      PE_gttx_nack,           // Recieved cmd was NACK'd

    // PHY Config Interface
    input                         PC_scram_disable,       // Scrambler Disable

    // OPLM Internal Signals
    input                         PPI_port_initialized,   // Link is init.
    input                         PPR_idle_selected,      // IDLE sequence selected (bind only)
    input                         PPR_idle2_selected,     // IDLE2 selected
    input                         PPI_mode_1x,            // Mode 1x Selected
    input       [LINK_WIDTH-1:0]  PPI_lane_sync           // Lanes Sync'd
    // }}} end port declarations ------------
  );

  // {{{ Localparams ------------------------
  // SRIO Protocol Parameters
  // ---------------------------
  localparam K_CHAR = 8'hBC; 
  localparam A_CHAR = 8'hFB; 
  localparam R_CHAR = 8'hFD;
  localparam M_CHAR = 8'h3C;
  localparam D0_0   = 8'h00;
  
  //Parameters for the CS Field Encodings (table 4-8 of PHY spec)
  localparam ENCODE_0_0  = 8'h67;  //D7.3  character
  localparam ENCODE_0_1  = 8'h78;  //D24.3 character
  localparam ENCODE_1_0  = 8'h7E;  //D30.3 character
  localparam ENCODE_1_1  = 8'hF8;  //D24.7 character

  //Parameters for the CS Field Marker of the IDLE2 Sequence
  localparam D21_5  = 8'hB5;  
  localparam D0_2   = 8'h40;  //Lane 0, LINK_WIDTH=4, !mode_1x
  localparam D1_2   = 8'h41;  //Lane 1, LINK_WIDTH=4, !mode_1x
  localparam D2_2   = 8'h42;  //Lane 2, LINK_WIDTH=4, !mode_1x
  localparam D3_2   = 8'h43;  //Lane 3, LINK_WIDTH=4, !mode_1x
  localparam D0_7   = 8'hE0;  //Lane 0, LINK_WIDTH=4, mode_1x
  localparam D1_7   = 8'hE1;  //Lane 1, LINK_WIDTH=4, mode_1x
  localparam D2_7   = 8'hE2;  //Lane 2, LINK_WIDTH=4, mode_1x
  localparam D3_7   = 8'hE3;  //Lane 3, LINK_WIDTH=4, mode_1x
  localparam D0_1   = 8'h20;  //Lane 0, LINK_WIDTH=2, !mode_1x
  localparam D1_1   = 8'h21;  //Lane 1, LINK_WIDTH=2, !mode_1x
  localparam D0_6   = 8'hC0;  //Lane 0, LINK_WIDTH=2, mode_1x
  localparam D1_6   = 8'hC1;  //Lane 1, LINK_WIDTH=2, mode_1x

  // OPLM TX Defined Parameters
  // ----------------------------
  localparam DATA_WIDTH_SYNC    = (LINK_WIDTH == 4) ? 128 : (LINK_WIDTH == 2) ? 64 : 32;
  localparam CHARIS_WIDTH_SYNC  = DATA_WIDTH_SYNC/8;
  localparam VALID_WIDTH        = (LINK_WIDTH == 4) ? 4   : (LINK_WIDTH == 2) ? 2  : 1;
  localparam VALID_DIVISOR      = (LINK_WIDTH == 4) ? 1   : (LINK_WIDTH == 2) ? 2  : 4;
  localparam VALID_HIGHBIT      = (LINK_WIDTH == 4) ? 3   : (LINK_WIDTH == 2) ? 1  : 0;

  // For idle the length of a synchronization seque is 5 cycles
  localparam SYNC_BYTES         = 20;
  localparam SYNC_CYCLES        = SYNC_BYTES/GT_BYTES;// 5 cycles to transmit
  localparam IDLE1_CCOMP_CYCLES = 1;                  // 1 cycles to transmit in IDLE1
  localparam IDLE2_CCOMP_CYCLES = 3;                  // 3 cycles to transmit in IDLE2
  localparam CSF_BYTES          = 40;                 // Bytes in the CS Field Total
  localparam CSF_CYCLES         = CSF_BYTES/GT_BYTES; // 40 characters, GT_BYTES characters/cycle
  localparam CSM_BYTES          = 8;                  // Bytes in the CS Field Marker only
  localparam CSM_CYCLES         = CSM_BYTES/GT_BYTES; 
  localparam CCOMP_WIDTH        = 11;                 // 11-bits is 1024
  localparam RAND_DF_MAX_CYCLES = 512/GT_BYTES;       // 128 cycles to transmit 512 D0.0s
  // }}} ------------------------------------

  // {{{ Wire Declarations ------------------
  // Clock Domain Crossing
  reg                           phy_rise_edge_det;
  reg                           phy_rise_edge_det_q;
  reg                           byte_idx;
  reg [DATA_WIDTH_SYNC-1:0]     tx_data_sync;
  reg [CHARIS_WIDTH_SYNC-1:0]   tx_charisk_sync;
  reg [VALID_WIDTH-1:0]         tx_valid_sync;

  reg [63:0]                    pt_tx_data_q;
  reg [7:0]                     pt_tx_charisk_q;
  reg [1:0]                     pt_tx_valid_q;
  reg                           pt_send_lreq_q = 0;
  reg                           pt_early_lreq_q = 0;

  reg                           ccomp_grant_sync;
  reg                           ccomp_req;
  reg                           lreq_sent;
  reg                           indicate_lreq_sent;
  wire                          lreq_complete;
  wire                          indicate_lreq_complete;
  reg   [2:0]                   sync_seq_ctr;

  // Striping Logic
  wire  [GT_BYTES*8-1:0]        stripe_d        [LINK_WIDTH-1:0];
  wire  [GT_BYTES-1:0]          stripe_isk_d    [LINK_WIDTH-1:0];
  wire  [GT_BYTES-1:0]          stripe_valid_d;
  reg   [GT_BYTES*8-1:0]        stripe          [LINK_WIDTH-1:0];
  reg   [GT_BYTES-1:0]          stripe_isk      [LINK_WIDTH-1:0];
  reg   [GT_BYTES-1:0]          stripe_valid;
  reg                           phy_is_valid;
  wire                          phy_is_valid_d;

  // Data Selection
  reg   [(GT_BYTES*8)-1:0]      lane_d          [LINK_WIDTH-1:0];
  reg   [GT_BYTES-1:0]          lane_isk        [LINK_WIDTH-1:0];
  reg   [GT_BYTES-1:0]          lane_valid      [LINK_WIDTH-1:0];
  reg   [(GT_BYTES*8)-1:0]      scram           [LINK_WIDTH-1:0];
  reg   [GT_BYTES-1:0]          scram_isk       [LINK_WIDTH-1:0];

  // Shared IDLE logic
  reg   [6:0]                   rng_curr;
  reg   [6:0]                   rng_next;
  reg   [2:0]                   a_m_ctr;
  wire                          a_m_ctr_eq0;
  wire                          a_m_load;
  wire  [GT_BYTES-1:0]          start_idle;

  // Clk Comp Logic
  wire                          ccomp_freq_ctr_max;
  reg   [CCOMP_WIDTH-1:0]       ccomp_freq_ctr;
  reg   [3:0]                   ccomp_ctr;
  reg                           send_ccomp;
  wire  [1:0]                   ccomp_cycles;

  // IDLE sequences
  reg   [(GT_BYTES*8)-1:0]      idle1;
  reg   [GT_BYTES-1:0]          idle1_isk;
  reg   [(GT_BYTES*8)-1:0]      idle2           [LINK_WIDTH-1:0];
  reg   [GT_BYTES-1:0]          idle2_isk       [LINK_WIDTH-1:0];
  wire  [(GT_BYTES*8)-1:0]      idle            [LINK_WIDTH-1:0];
  wire  [GT_BYTES-1:0]          idle_isk        [LINK_WIDTH-1:0];
  reg                           cs_field;
  reg                           cs_field_start;
  reg                           cs_field_q;
  reg                           send_sync;
  reg                           valid_send_lreq;
  reg                           shift_sync_seq;
  reg   [7:0]                   rand_df_ctr;
  wire                          mask_idles;
  wire                          send_csfm;
  wire                          send_csf;
  reg                           send_lreq_sync;
  reg                           early_lreq_sync;
  reg                           send_lreq_sync_q;
  wire  [GT_BYTES*8-1:0]        sync_seq;
  wire  [GT_BYTES-1:0]          sync_seq_isk;

  // Output
  reg                           tx_idle2_selected;
  reg                           tx_idle2_selected_q;
  wire  [DATA_WIDTH-1:0]        gttx_data_d;
  wire  [CHARIS_WIDTH-1:0]      gttx_charisk_d;
  // }}} -------------------------------------

  // {{{ Clock Domain Crossing --------------
  //phy_clk rising edge detect circuit used to reset the byte_idx counter
  //The phy_rise_edge_det signal samples toggles in the phy_clk domain,
  //The phy_rise_edge_det_q signal is sampled in the gt_pcs_clk domain in order to
  //detect the edge change in the gt_pcs_clk domain. These to signals in
  //conjunction detect the rising edge of every phy_clk cycle to reset
  //the byte index we are sampling from out of the tx_data bus and
  //corresponding sideband signals.  This is used to determine loading 
  //conditions for the byte_idx ctr because each domain can be reset
  //independently.
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      phy_rise_edge_det <= #TCQ 1'b0;
    end else begin
      phy_rise_edge_det <= #TCQ ~phy_rise_edge_det;
    end
  end

  //Start out with 1 so the byte_idx will immediately load after a reset
  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      phy_rise_edge_det_q  <= #TCQ 1'b1;
    end else begin
      phy_rise_edge_det_q  <= #TCQ phy_rise_edge_det;
    end
  end

  wire byte_idx_load = phy_rise_edge_det_q != phy_rise_edge_det;

  // Based on the link width increment through the byte locations
  // of the data in the phy clock domain. This is only needed for x1
  // cores where the gt_pcs_clk is faster than phy_clk. Because the edge 
  // detector will not be able to detect the rising edge until a cycle later, 
  // the load value of the byte counter will need to start at the second 
  // half of the dword.
  // when the sync sequence is being sent, the lreq needs to hold at byte 1
  // to send the link request aligned in the proper order
  always @(posedge gt_pcs_clk) begin
    if (byte_idx_load) begin
      byte_idx <= #TCQ (send_sync) ? ~sync_seq_ctr[0] : 0;
    end else begin
      byte_idx <= #TCQ ~byte_idx;
    end
  end

  // Based on the link width create the logic to cross domains
  generate if (LINK_WIDTH == 1) begin: x1_sync_gen
    // gt_pcs_clk*2 == phy_clk
    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        // Only need a reset of the control bits
        tx_valid_sync        <= #TCQ 0;
      end else begin
        tx_data_sync         <= #TCQ PT_tx_data[(byte_idx*32)+:32];
        tx_charisk_sync      <= #TCQ PT_tx_charisk[(byte_idx*4)+:4];
        tx_valid_sync        <= #TCQ PT_tx_valid[byte_idx];
      end
    end

  end else if (LINK_WIDTH == 2) begin: x2_sync_gen
    // gt_pcs_clk == phy_clk
    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        // Only need a reset of the control bits
        tx_valid_sync        <= #TCQ 0;
      end else if (PPI_mode_1x) begin
        tx_data_sync         <= #TCQ PT_tx_data[(byte_idx*32)+:32];
        tx_charisk_sync      <= #TCQ PT_tx_charisk[(byte_idx*4)+:4];
        tx_valid_sync        <= #TCQ PT_tx_valid[byte_idx];
      end else begin
        tx_data_sync          <= #TCQ PT_tx_data;
        tx_charisk_sync       <= #TCQ PT_tx_charisk;
        tx_valid_sync         <= #TCQ PT_tx_valid;
      end
    end
  end else if (LINK_WIDTH == 4) begin: x4_sync_gen
    // gt_pcs_clk/2 == phy_clk
    always @(posedge phy_clk) begin
      if (phy_rst_q) begin
        // Only need a reset of the control bits
        pt_tx_valid_q      <= #TCQ 0;
        pt_send_lreq_q     <= #TCQ 0;
        pt_early_lreq_q    <= #TCQ 0;
      end else begin
        pt_tx_data_q       <= #TCQ PT_tx_data;
        pt_tx_charisk_q    <= #TCQ PT_tx_charisk;
        pt_tx_valid_q      <= #TCQ PT_tx_valid;
        pt_send_lreq_q     <= #TCQ PT_send_lreq;
        pt_early_lreq_q    <= #TCQ PT_tx_early_lreq;
      end
    end

    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        // Only need a reset of the control bits
        tx_valid_sync        <= #TCQ 0;
      end else if (PPI_mode_1x) begin
        tx_data_sync         <= #TCQ PT_tx_data[(byte_idx*32)+:32];
        tx_charisk_sync      <= #TCQ PT_tx_charisk[(byte_idx*4)+:4];
        tx_valid_sync        <= #TCQ PT_tx_valid[byte_idx];
      end else begin
        tx_data_sync         <= #TCQ {pt_tx_data_q,    PT_tx_data};
        tx_charisk_sync      <= #TCQ {pt_tx_charisk_q, PT_tx_charisk};
        tx_valid_sync        <= #TCQ (!pt_send_lreq_q && PT_send_lreq) ? 
                                        {pt_tx_valid_q, 2'b00} :
                                        {pt_tx_valid_q, PT_tx_valid};
      end
    end
  end endgenerate

  //Synchronize Incoming signals to the GT Clock
  always @(posedge gt_pcs_clk) begin    
    if (gt_pcs_rst_q) begin
      ccomp_grant_sync <= #TCQ 0;
      send_lreq_sync   <= #TCQ 0;
      early_lreq_sync  <= #TCQ 0;
    end else begin
      ccomp_grant_sync <= #TCQ PT_ccomp_grant;

      if (!PPI_mode_1x && LINK_WIDTH == 4) begin
        send_lreq_sync  <= #TCQ pt_send_lreq_q;
        early_lreq_sync <= #TCQ pt_early_lreq_q;
      end else begin
        send_lreq_sync  <= #TCQ PT_send_lreq;
        early_lreq_sync <= #TCQ PT_tx_early_lreq;
      end
    end
  end

  //Synchronize the Outgoing signals to the PHY clock
  always @(posedge phy_clk) begin    
    if (phy_rst_q) begin
      PPT_ccomp_req <= #TCQ 0;
      PPT_lreq_sent <= #TCQ 0;
    end else begin
      PPT_ccomp_req <= #TCQ ccomp_req;
      PPT_lreq_sent <= #TCQ indicate_lreq_sent;
    end
  end  
  // }}} end Clock Domain Crossing ----------

  // {{{ Lane Striping ----------------------
  // Stripe the incoming data across all active lanes
  // Generate the striping logic for each lane based on the link width
  genvar std_ii; // striping _d 
  genvar stb_ii; // striping bytes
  generate for (stb_ii=0; stb_ii < GT_BYTES; stb_ii=stb_ii+1) begin: stripe_d_byte_gen
    for (std_ii=0; std_ii < LINK_WIDTH; std_ii=std_ii+1) begin: stripe_d_lane_gen
      assign stripe_d[(LINK_WIDTH-1)-std_ii][(stb_ii*8)+:8] = tx_data_sync[((LINK_WIDTH*8*stb_ii)+(std_ii*8))+:8];
      assign stripe_isk_d[(LINK_WIDTH-1)-std_ii][stb_ii]    = tx_charisk_sync[LINK_WIDTH*stb_ii+std_ii];
    end //end for (stb_ii < GT_BYTES)

    assign stripe_valid_d[stb_ii] = (phy_is_valid) ? 1'b0 : tx_valid_sync[stb_ii/VALID_DIVISOR];
  end endgenerate// end for (std_ii < LINK_WIDTH)
    
  genvar st_ii; // striping
  generate for (st_ii=0; st_ii < LINK_WIDTH; st_ii=st_ii+1) begin: stripe_gen
    always @(posedge gt_pcs_clk) begin
      // No need to reset the data bits
      if (PPI_mode_1x) begin
        stripe[st_ii]        <= #TCQ tx_data_sync[31:0];
        stripe_isk[st_ii]    <= #TCQ tx_charisk_sync[3:0];
      end else begin
        stripe[st_ii]        <= #TCQ stripe_d[st_ii];
        stripe_isk[st_ii]    <= #TCQ stripe_isk_d[st_ii];
      end
    end
  end endgenerate //end for (st_ii < LINK_WIDTH)
  
  wire mask_last_lreq = (indicate_lreq_sent && !early_lreq_sync && PPI_mode_1x && (sync_seq_ctr < 4));

  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      stripe_valid  <= #TCQ 0;
    end else begin
      // If there is a link request to send, once the link request is sent 
      // clear the valid bus until the handshake is complete and new data is 
      // present to avoid sending two of the same link request
      if (((lreq_complete || lreq_sent) || mask_last_lreq) && send_lreq_sync) begin
        stripe_valid <= #TCQ 0;

      end else if (PPI_mode_1x) begin
        stripe_valid <= #TCQ {GT_BYTES{tx_valid_sync[0]}};

      // In x4 mode two long control symbol can fit on one cycle which means when
      // a link request needs to be sent then the lreq can be sent twice since it
      // will be striped while the SYNC seq is being sent. To avoid this, mask 
      // off the lower two bits of the valid data
      end else if ((send_lreq_sync) && (LINK_WIDTH == 4)) begin
        stripe_valid <= #TCQ (!shift_sync_seq) ? 4'b1100 : 4'b0011;

      end else begin
        stripe_valid <= #TCQ stripe_valid_d;
      end
    end
  end
  
  //Evaluation Core Logic
  //Only generate this is EVAL is set.  This will mask off the incoming valid
  //to be always 0 so no data will be sent out only idles.
  generate if (EVAL) begin : validlogic_gen
    //The eval logic can not be reset
    srio_gen2_v4_1_16_eval_gt_pcs_clk  #(
      .TCQ (TCQ),
      .MODE_XG (MODE_XG)
    ) valid_inst (
      .flag (phy_is_valid_d),
      .rst  (1'b0),
      .clk  (gt_pcs_clk)
     );
  end else begin: passthrough_gen
    assign phy_is_valid_d = 0;
  end endgenerate
  always @(posedge gt_pcs_clk) begin
    phy_is_valid <= #TCQ phy_is_valid_d;
  end

  //*COVERPOINT
  //(cp_stripe_valid):Valid Data arrives on byte 0, both bytes, and no bytes, data arriving from the 
  // ollm tx on byte 1 only is invalid
  // }}} Lane Striping ----------------------
  
  // {{{ + Idle Sequence Generator + ------------
  // Save the PP_idle2_selected signal.  When important functions are being
  // performed. This needs to remain stable for the idle sequence generation
  // to remain spec compliant
  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      tx_idle2_selected   <= #TCQ IDLE2;
      tx_idle2_selected_q <= #TCQ IDLE2;
    end else begin
      if (!send_ccomp) begin
        tx_idle2_selected <= #TCQ PPR_idle2_selected;
      end
      tx_idle2_selected_q <= #TCQ tx_idle2_selected;
    end
  end

  //*COVERAGE*
  //(cp_idle2_changes_during_ccomp): See a change in the idle mode while a clock comp is being sent
  // for the last idle mode
  
  //Linear Feedback Shift Register (LFSR)
  //Shift to the next state according to the function f(x) = x^7 ^ x^6 + 1
  //the following values of rng_next is based on a two bit parallelzation 
  //of f(x).  This polynomail is take directly from the PHY layer spec.
  //See the Idle1 sequence section for more details.  
  //rng = random number generator
  always @(*) begin
    rng_next[0] = rng_curr[6] ^ rng_curr[2];
    rng_next[1] = rng_curr[5] ^ rng_curr[1];
    rng_next[2] = rng_curr[1];
    rng_next[3] = rng_curr[2];
    rng_next[4] = rng_curr[3];
    rng_next[5] = rng_curr[4];
    rng_next[6] = rng_curr[5];
  end

  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      rng_curr <= #TCQ -1; //initialize to all 1's
    end else begin
      rng_curr <= #TCQ rng_next;
    end
  end

  //Down-Counter for placement of A or M special characters
  //If we are starting an IDLE sequence we cant start with a special
  //character, this is specific to idle2 but can be used for both IDLE
  //sequences
  assign a_m_ctr_eq0 = (a_m_ctr == 0) && !(|start_idle);

  // When loading the a_m_ctr in IDLE2 there is the additional requirements of:
  // 1. The random data field starts over after the Command and Status Field
  // 2. The random data field starts over after a clock compensation sequence.
  // 3. A sync sequence doesnt need to be sent
  wire   a_m_load_any_idle = a_m_ctr_eq0 || |start_idle;
  wire   a_m_load_idle2    = a_m_load_any_idle || cs_field || send_ccomp || 
                             (send_lreq_sync && !lreq_sent && |stripe_valid);
  assign a_m_load          = tx_idle2_selected ? a_m_load_idle2 : a_m_load_any_idle;
  
  //*ASSERTION*
  // (ap_a_m_underflow): a_m_ctr does not underflow
  // (ap_a_m_overcount): a_m_ctr does not go above the max value, 6

  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      a_m_ctr <= #TCQ -1; //Initialize to all 1's

    end else begin
      // Load with a new random value of 5 or 4. These numbers were chosen
      // to be sure there are at least 16-31 characters between A's for a 4 byte
      // GT interface.
      if (a_m_load)
        a_m_ctr <= #TCQ {1'b1, 1'b0, (rng_curr[4])};
      else  
        a_m_ctr <= #TCQ a_m_ctr - 1'b1;
    end
  end

  //clock compensation sequence frequency of events counter
  assign ccomp_freq_ctr_max = ccomp_freq_ctr[CCOMP_WIDTH-1];

  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      ccomp_freq_ctr <= #TCQ 0;
    end else begin 
      if (ccomp_freq_ctr_max) begin
        ccomp_freq_ctr <= #TCQ 0; 
      end else begin
        ccomp_freq_ctr <= #TCQ ccomp_freq_ctr + 1'b1;
      end
    end
  end
  
  // Select the appropriate number of cycles to transmit the clk comp
  // sequence depending on the idle mode.
  assign ccomp_cycles = (tx_idle2_selected) ? IDLE2_CCOMP_CYCLES-1 : 
                                              IDLE1_CCOMP_CYCLES-1;

  // Start sending the clk comp when we know there will not a be an A required
  // If there was a K character on the idle it was from the a_m_ctr_eq0 being
  // valid just before the ccomp grant arrived, so wait a cycle to maintain
  // the requirement that it must have 4 D0 characters following.

  // Before sending the ccomp sequence we need to meet the following criteria:
  // 1. There has to be enough D0 characters before the ccomp starts, 4 cycles 
  // will be 16 which is the min req.
  wire start_ccomp_seq = ccomp_req && ccomp_grant_sync && (a_m_ctr > 3);
  
  //*ASSERTION*
  //(ap_ccomp_grant_only_with_req): If the clk comp is granted then there must be a request

  //*COVERAGE*
  //(cp_ccomp_a_m_ctr_1, cp_ccomp_a_m_ctr_0): See a ccomp request that is granted when 
  // the a_m_ctr is 1 and 0, and loading

  //*COVERAGE*
  //(cp_ccomp_csf_starts): See a ccomp request that is granted when the csf field
  // starts

  //(cp_ccomp_csf_enbd): See a ccomp request that is granted when the csf field
  // ends

  // Only count ccomp cycles in IDLE2 mode, in IDLE1 it only takes one cycle to send
  // the ccomp sequence.
  wire ccomp_ctr_rst;

  generate if (IDLE2) begin: ccomp_ctr_gen
    assign ccomp_ctr_rst = (ccomp_ctr == ccomp_cycles);

    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        send_ccomp <= #TCQ 0;
      end else begin
        if (ccomp_ctr_rst) begin
          send_ccomp <= #TCQ 1'b0;

        end else if (start_ccomp_seq) begin
          send_ccomp <= #TCQ 1'b1;
        end
      end
    end

    //count the number of cycles of clock comp sent
    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        ccomp_ctr <= #TCQ 0;
      end else begin
        if (ccomp_ctr_rst)
          ccomp_ctr <= #TCQ 0;
        else if (send_ccomp)
          ccomp_ctr <= #TCQ ccomp_ctr + 1'b1;
      end
    end
  
  end else begin: no_ccomp_ctr_gen
    // Tie off globally used signals created in this block
    always @(posedge gt_pcs_clk) begin
      send_ccomp <= #TCQ 0;
    end
    assign ccomp_ctr_rst = 0;
  end endgenerate
  
  //*ASSERTION*
  //(ap_ccomp_underflow): Clock Compensation Cycle counter does not underflow
  //(ap_ccomp_overflow): Clock Compensation Cycle counter does not overflow

  // Tweak when ccomp_req is deasserted in order to get data through the pipe
  // quickly by subtracting cycles for latency. In idle1 mode since the ccomp
  // is only two cycles we can deassert the request as soon as it is granted.
  wire deassert_ccomp_req = tx_idle2_selected ? send_ccomp : 
                                                start_ccomp_seq;

  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      ccomp_req <= #TCQ 0;
    end else begin
      if (deassert_ccomp_req) begin
        ccomp_req <= #TCQ 0;
      end else if (ccomp_freq_ctr_max) begin
        ccomp_req <= #TCQ 1;
      end
    end
  end
  //*ASSERTION*
  //(ap_ccomp_asserts_within_5000): with divided counter set the ccomp request must
  // assert after every 4096 characters

  //*ASSERTION*
  //(ap_ccomp_asserts_too_frequently): a ccomp request should not bee seen less than
  // the designated amount of time

  //*ASSERTION*
  //(ap_ccomp_granted_ontime): After a clock compensation request, it must be granted within 904 
  // characters.

  //*COVERAGE*
  // (cp_start_idle): An idle sequence starts on each bytes on a lane
  // Any other combination of this signal is invalid

  // Determine if there is a start of a idle sequence on the next dword.
  assign start_idle[0] = stripe_valid_d[1] && !stripe_valid_d[0] && !send_lreq_sync_q;
  assign start_idle[1] = stripe_valid_d[2] && !stripe_valid_d[1] && !send_lreq_sync_q;
  assign start_idle[2] = stripe_valid_d[3] && !stripe_valid_d[2] && !send_lreq_sync_q;
  assign start_idle[3] = stripe_valid[0]   && !stripe_valid_d[3] && !send_lreq_sync_q;
  
  // {{{ IDLE1 Sequence Generator
  //Declare those wires used only for the IDLE1 sequence generator.
  //These are created outside the scope of the generate in order to assist
  //in coverage in the bind files.  This enables automatic binding and
  //eliminates the need for heirarchical references.
  wire [GT_BYTES-1:0] i1_send_k;
  wire [GT_BYTES-1:0] i1_send_a;
  wire [GT_BYTES-1:0] i1_send_r;

  //If IDLE1 mode is supported, generate the logic that generates IDLE1
  //sequences.
  genvar i1r_ii; // i1_rand_* 
  generate if (IDLE1) begin: idle1_seq_gen
    reg [(GT_BYTES*8)-1:0]  i1_rand;

    //The clock comp seq is written so the LSB is selected first
    wire [31:0] IDLE1_CCOMP_SEQ = {K_CHAR, R_CHAR, R_CHAR, R_CHAR}; 

    // Use bits in the lfsr to randomly select which character to send on
    // which bit.  If there is an A to be sent, that is always selected over
    // a K or R. A K must be selected if it is the start of the IDLE1 sequence.
    // The A is randomly placed on a byte. The rng indexes selected are
    // completely random and can easily be replaced with any bits
    assign i1_send_k[0]  = (!i1_send_a[0] && rng_curr[2]) || start_idle[0];
    assign i1_send_k[1]  = (!i1_send_a[1] && rng_curr[0]) || start_idle[1];
    assign i1_send_k[2]  = (!i1_send_a[2] && rng_curr[6]) || start_idle[2];
    assign i1_send_k[3]  = (!i1_send_a[3] && rng_curr[4]) || start_idle[3];

    assign i1_send_r[0]  = !i1_send_a[0] && !rng_curr[2] && !start_idle[0];
    assign i1_send_r[1]  = !i1_send_a[1] && !rng_curr[0] && !start_idle[1];
    assign i1_send_r[2]  = !i1_send_a[2] && !rng_curr[6] && !start_idle[2];
    assign i1_send_r[3]  = !i1_send_a[3] && !rng_curr[4] && !start_idle[3];

    assign i1_send_a[0]  = a_m_ctr_eq0 && (!rng_curr[1] && !rng_curr[3]) && !start_idle[0];
    assign i1_send_a[1]  = a_m_ctr_eq0 && (!rng_curr[1] && rng_curr[3])  && !start_idle[1];
    assign i1_send_a[2]  = a_m_ctr_eq0 && (rng_curr[1] && !rng_curr[3])  && !start_idle[2];
    assign i1_send_a[3]  = a_m_ctr_eq0 && (rng_curr[1] && rng_curr[3])   && !start_idle[3];

    //*ASSERTION*   
    //(ap_i1_onehot): When selecting K, As, and Rs, only one send_* indicator can be
    // asserted for each byte

    // Populate the i1_rand bus for the idle field's 4 bytes
    for (i1r_ii = 0; i1r_ii< GT_BYTES; i1r_ii=i1r_ii+1) begin: i1_rand_gen
      always @(*) begin
        case ({i1_send_k[i1r_ii],i1_send_a[i1r_ii],i1_send_r[i1r_ii]})
          3'b100: i1_rand[i1r_ii*8+:8] = K_CHAR;
          3'b010: i1_rand[i1r_ii*8+:8] = A_CHAR;
          3'b001: i1_rand[i1r_ii*8+:8] = R_CHAR;
          default:i1_rand[i1r_ii*8+:8] = 8'bX;
        endcase
      end
    end

    // Select the clock comp sequence or the random idle sequence.
    // Only keep track of one lane since all should be transmitted identically
    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        idle1     <= #TCQ {K_CHAR, i1_rand[23:0]};
        idle1_isk <= #TCQ {GT_BYTES{1'b1}};
      end else begin
        idle1     <= #TCQ (start_ccomp_seq) ? IDLE1_CCOMP_SEQ : i1_rand;
        idle1_isk <= #TCQ {GT_BYTES{1'b1}};
      end
    end

  end //end if (IDLE1)
  else begin: no_idle1_seq_gen
    //Tie off these wires for the bind files.
    assign i1_send_k = 0;
    assign i1_send_a = 0;
    assign i1_send_r = 0;
  end endgenerate
  // }}} IDLE1 Sequence Generator
  
  // {{{ IDLE2 Sequence Generator
  //Declare those wires used only for the IDLE2 sequence generator.
  //These are created outside the scope of the generate in order to assist
  //in coverage in the bind files.  This enables automatic binding and
  //eliminates the need for heirarchical references.
  wire  [GT_BYTES-1:0]      i2_send_a;
  wire  [GT_BYTES-1:0]      i2_send_m;
  reg   [GT_BYTES-1:0]      csf_ctr;
  reg   [(GT_BYTES*8)-1:0]  i2_rand;
  reg   [GT_BYTES-1:0]      i2_isk_rand;
  wire  [GT_BYTES*8-1:0]    csf_select_encoded [LINK_WIDTH-1:0];
  wire  [LINK_WIDTH-1:0]    send_ack;
  wire  [LINK_WIDTH-1:0]    send_nack;
  wire  [LINK_WIDTH-1:0]    send_cmd;
  reg   [LINK_WIDTH-1:0]    ack_pending;
  reg   [LINK_WIDTH-1:0]    nack_pending;
  reg   [LINK_WIDTH-1:0]    cmd_pending;
  
  genvar cs_ii;  // cs field
  genvar i2_ii;  // idle2 gen
  genvar i2r_ii; // i2_rand_* gen
  //If IDLE2 mode is supported, generate the logic used to generate the IDLE2
  //sequence.
  generate 
    if (IDLE2) begin: idle2_seq_gen
      wire          rand_df_reset;
      reg           idle_frame_toggle;
      wire  [63:0]  csfm              [LINK_WIDTH-1:0];
      wire  [7:0]   csfm_isk;
      reg   [31:0]  csfield           [LINK_WIDTH-1:0];
      wire  [63:0]  tx_csf            [LINK_WIDTH-1:0];

      // {{{ CS Field Creation
      //M, D, D, D, D, D is added on the end of the cc seq. since a cc seq must
      //be followed by an idle frame which must start with an M and and idle
      //seq can not terminate with < 4 D's following an M.
      wire [95:0] IDLE2_CCOMP_SEQ = {K_CHAR, R_CHAR, R_CHAR, R_CHAR,
                                     M_CHAR, D0_0,   D0_0,   D0_0, 
                                     D0_0,   D0_0,   D0_0,   D0_0};

      wire [11:0] IDLE2_CCOMP_SEQ_ISK = {5'b11111, 7'b0000000};

      for (cs_ii = 0; cs_ii < LINK_WIDTH; cs_ii=cs_ii+1) begin: csf_gen
        //Whenever a ack/nack is detected latch it until it is sent
        reg [1:0] tap_m1_cmd;
        reg [1:0] tap_p1_cmd;
        reg       reset_emphasis;
        reg       preset_emphasis;

        // Look for the rising edge of an ack/nack to know when to send one in
        // the next cs_field
        assign send_ack[cs_ii]   = !ack_pending[cs_ii] && PE_gttx_ack[cs_ii];
        assign send_nack[cs_ii]  = !nack_pending[cs_ii] && PE_gttx_nack[cs_ii];
        assign send_cmd[cs_ii]   = !cmd_pending[cs_ii] && PE_gttx_cmd[cs_ii];
      
        //*COVERAGE*
        //(cp_send_ack): Send an Ack in the command and status field
        //(cp_send_nack): Send an Nack in the command and status field
        //(cp_send_cmd): Send a command in the command and status field
        
        //*ASSERTION*
        //(ap_send_idle2_only): A send command can only occur in idle2 mode

       //*ASSERTION*
       //(ap_ack_deasserts, ap_nack_deasserts, ap_cmd_deasserts): 
       // A pending command for the cs field can only drop once a csfield is sent

        // An ack/nack is sent when beat 
        wire resp_sent = send_csf && (csf_ctr == CSF_CYCLES-1); //last beat of the CSF

        // Set and ack on the rising edge of PE_gttx_ack, release it when that
        // beat of the CSF is sent.
        always @(posedge gt_pcs_clk) begin
          if (gt_pcs_rst_q) begin
            ack_pending[cs_ii] <= #TCQ 0;
          end else begin
            if (resp_sent) begin
              ack_pending[cs_ii] <= #TCQ 0;
            end else if (send_ack[cs_ii]) begin
              ack_pending[cs_ii] <= #TCQ 1;
            end
          end
        end

        // Set and nack on the rising edge of PE_gttx_ack, release it when that
        // beat of the CSF is sent.
        always @(posedge gt_pcs_clk) begin
          if (gt_pcs_rst_q) begin
            nack_pending[cs_ii] <= #TCQ 0;
          end else begin
            if (resp_sent) begin
              nack_pending[cs_ii] <= #TCQ 0;
            end else if (send_nack[cs_ii]) begin
              nack_pending[cs_ii] <= #TCQ 1;
            end
          end
        end

        // Register a command to send and hold it till a CSF is sent
        always @(posedge gt_pcs_clk) begin
          if (gt_pcs_rst_q) begin
            cmd_pending[cs_ii]  <= #TCQ 0;
            tap_m1_cmd          <= #TCQ 0;
            tap_p1_cmd          <= #TCQ 0;
            preset_emphasis     <= #TCQ 0;
            reset_emphasis      <= #TCQ 0;
          end else begin
            if (resp_sent) begin
              cmd_pending[cs_ii]  <= #TCQ 0;
              tap_m1_cmd          <= #TCQ 0;
              tap_p1_cmd          <= #TCQ 0;
              preset_emphasis     <= #TCQ 0;
              reset_emphasis      <= #TCQ 0;

            end else if (send_cmd[cs_ii]) begin
              cmd_pending[cs_ii]  <= #TCQ PE_gttx_cmd[cs_ii];
              tap_m1_cmd          <= #TCQ PE_gttx_tap_m1_cmd[cs_ii*2+:2];
              tap_p1_cmd          <= #TCQ PE_gttx_tap_p1_cmd[cs_ii*2+:2];
              preset_emphasis     <= #TCQ PE_gttx_preset_emphasis[cs_ii];
              reset_emphasis      <= #TCQ PE_gttx_preset_emphasis[cs_ii];
            end
          end
        end
        
        // Only update these bits if we are not currently transmitting the
        // cs_field, otherwise the bitwise complement will be corrupt.
        // It does not need a reset since it will all be valid by the first
        // time it is transmitted and all the signals which populate this
        // field have a reset
        always @(posedge gt_pcs_clk) begin
          if (!cs_field) begin
            csfield[cs_ii][31]    <= #TCQ cmd_pending[cs_ii];                //Command Present
            csfield[cs_ii][30]    <= #TCQ 1'b0;                              //Implementation Defined
            csfield[cs_ii][29]    <= #TCQ &PPI_lane_sync;                    //Receiver is Trained
            csfield[cs_ii][28]    <= #TCQ !PC_scram_disable;                 //Scrambling Enabled
            csfield[cs_ii][27:26] <= #TCQ PE_gttx_tap_m1_status[cs_ii*2+:2]; //Tap (-1) Status
            csfield[cs_ii][25:24] <= #TCQ PE_gttx_tap_p1_status[cs_ii*2+:2]; //Tap (+1) Status
            csfield[cs_ii][23:8]  <= #TCQ 16'h00;                            //Reserved
            csfield[cs_ii][7:6]   <= #TCQ tap_m1_cmd;                        //Tap (-1) 
            csfield[cs_ii][5:4]   <= #TCQ tap_p1_cmd;                        //Tap (+1)
            csfield[cs_ii][3]     <= #TCQ reset_emphasis;                    //Reset Emphasis
            csfield[cs_ii][2]     <= #TCQ preset_emphasis;                   //Preset Emphasis
            csfield[cs_ii][1]     <= #TCQ ack_pending[cs_ii];                //Ack
            csfield[cs_ii][0]     <= #TCQ nack_pending[cs_ii];               //Nack
          end
        end

        //Create the 64-bit CSF as indicated by the PHY Spec section 4.7.4.1.3
        //(Idle2 Command and Status Field)
        assign tx_csf[cs_ii] = {csfield[cs_ii], ~csfield[cs_ii]};
      end //end for
      // }}} end CS Field Creation

      // {{{ CSENCODE Function
      //the csencode function encodes the CS Field using 4 bits at a time to
      //create a 16-bit value as indicated by the PHY Spec in table 4-8
      function [31:0] csencode (
        input [7:0] x //value to encode
      );
        begin
          case(x[1:0])
            2'b00: csencode[7:0] = ENCODE_0_0;
            2'b01: csencode[7:0] = ENCODE_0_1;
            2'b10: csencode[7:0] = ENCODE_1_0;
            2'b11: csencode[7:0] = ENCODE_1_1;
          endcase
          case(x[3:2])
            2'b00: csencode[15:8] = ENCODE_0_0;
            2'b01: csencode[15:8] = ENCODE_0_1;
            2'b10: csencode[15:8] = ENCODE_1_0;
            2'b11: csencode[15:8] = ENCODE_1_1;
          endcase
          case(x[5:4])
            2'b00: csencode[23:16] = ENCODE_0_0;
            2'b01: csencode[23:16] = ENCODE_0_1;
            2'b10: csencode[23:16] = ENCODE_1_0;
            2'b11: csencode[23:16] = ENCODE_1_1;
          endcase
          case(x[7:6])
            2'b00: csencode[31:24] = ENCODE_0_0;
            2'b01: csencode[31:24] = ENCODE_0_1;
            2'b10: csencode[31:24] = ENCODE_1_0;
            2'b11: csencode[31:24] = ENCODE_1_1;
          endcase
        end
      endfunction
      // }}} CSENCODE Function

      // {{{ CSFM Definitions
      //generate the appropriate CS fields based on the lane width
      //the LSB goes out first and the MSB goes out last when selected
      if (LINK_WIDTH == 4) begin: idle2_x4_csf_gen
        //when the link width is 4x, and mode_1x is true,
        //lanes 1 and 3 are not transmitted on, so we do not need
        //to include the trained csfm for these lanes
        assign csfm[0] = (PPI_mode_1x) ? {M_CHAR, M_CHAR, M_CHAR, M_CHAR, 
                                          D21_5, D0_7, D21_5, ~D0_7} :
                                         {M_CHAR, M_CHAR, M_CHAR, M_CHAR,
                                          D21_5, D0_2, D21_5, ~D0_2};  
       
        assign csfm[1] = {M_CHAR, M_CHAR, M_CHAR, M_CHAR, 
                          D21_5, D1_2, D21_5, ~D1_2};

        assign csfm[2] = (PPI_mode_1x) ? {M_CHAR, M_CHAR, M_CHAR, M_CHAR,
                                          D21_5, D2_7, D21_5, ~D2_7} :
                                         {M_CHAR, M_CHAR, M_CHAR, M_CHAR,
                                          D21_5, D2_2, D21_5, ~D2_2}; 

        assign csfm[3] = {M_CHAR, M_CHAR, M_CHAR, M_CHAR,
                          D21_5, D3_2, D21_5, ~D3_2}; 

      end else if (LINK_WIDTH == 2) begin: idle2_x2_csf_gen
        assign csfm[0] = (PPI_mode_1x) ? {M_CHAR, M_CHAR, M_CHAR, M_CHAR,
                                          D21_5, D0_6, D21_5, ~D0_6} :
                                         {M_CHAR, M_CHAR, M_CHAR, M_CHAR,
                                          D21_5, D0_1, D21_5, ~D0_1};  

        assign csfm[1] = (PPI_mode_1x) ? {M_CHAR, M_CHAR, M_CHAR, M_CHAR,
                                          D21_5, D1_6, D21_5, ~D1_6} :
                                         {M_CHAR, M_CHAR, M_CHAR, M_CHAR,
                                          D21_5, D1_1, D21_5, ~D1_1};                                             
      end else if (LINK_WIDTH == 1) begin: idle2_x1_csf_gen
        assign csfm[0] = {M_CHAR, M_CHAR, M_CHAR, M_CHAR,
                          D21_5, D0_0, D21_5, ~D0_0};
      end
      // }}} CSFM Definitions

      //Mark only the M's in the CSFM as K character. This will be the same
      //across all command and status fields for each lane
      assign csfm_isk = 8'b1111_0000;

      // Determine when to mask off the idle sequence for termination based on
      // the operating link width. Since the clock frequency changes and no
      // matter what we need 4 D0.0 characters at the end of a idle we need to
      // check the incoming valid at different stages back in the pipe.
      wire mask_conditions = !send_ccomp && !cs_field_q && !cs_field;
      
      // Because a x4 core operates on 128 bytes of data, any combination of the
      // valid is possible. So in that case idles need to be masked on two cycles
      if (LINK_WIDTH == 4) begin: x4_mask_gen
        assign mask_idles = (!PPI_mode_1x) ? 
                              (mask_conditions && (|stripe_valid || |tx_valid_sync)) || 
                              (!send_ccomp && |stripe_valid) : 
                              (mask_conditions && tx_valid_sync);
      end else begin: other_mask_gen
        assign mask_idles = (mask_conditions && tx_valid_sync);
      end

      //Use random bits from the lfsr to select which byte to put an A/M on
      //this is only done when the down counter reaches 0
      //The bits from the RNG 6, and 1, and 5 are randomly selected, these could be
      //any bits, however between i2_send_*0's or i2_send_*1's they need to use
      //the same bits so no two are selected at once.
      assign i2_send_a[0] = a_m_ctr_eq0 && !rng_curr[6] && !rng_curr[1] && !rng_curr[5];
      assign i2_send_a[1] = a_m_ctr_eq0 && !rng_curr[6] && !rng_curr[1] &&  rng_curr[5];
      assign i2_send_a[2] = a_m_ctr_eq0 && !rng_curr[6] &&  rng_curr[1] && !rng_curr[5];
      assign i2_send_a[3] = a_m_ctr_eq0 && !rng_curr[6] &&  rng_curr[1] &&  rng_curr[5];

      assign i2_send_m[0] = a_m_ctr_eq0 && rng_curr[6] && !rng_curr[1] && !rng_curr[5]; 
      assign i2_send_m[1] = a_m_ctr_eq0 && rng_curr[6] && !rng_curr[1] &&  rng_curr[5]; 
      assign i2_send_m[2] = a_m_ctr_eq0 && rng_curr[6] &&  rng_curr[1] && !rng_curr[5]; 
      assign i2_send_m[3] = a_m_ctr_eq0 && rng_curr[6] &&  rng_curr[1] &&  rng_curr[5]; 

      //*ASSERTION*
      //(ap_i2_onehot): sending an A || M should never indicate to send both.

      //*COVERAGE*
      //(cp_i2_send_a_bytes): See an A need to be send on every byte
      //(cp_i2_send_m_bytes): See and M need to be sent on every byte

      //Create an idle frame toggle switch. This has a value of 1 when it
      //needs to transmit the random data field of the idle frame. This has
      //a value of 0 when it is transmitting the Command and Status Field
      //Rand data field transmission starts after valid data or after the cs
      //field is transmitted.
      //The CS field always starts after the random data field counter reaches
      //its max value of 128 indicating ~508 rand bytes have been sent.
      assign rand_df_reset = (|tx_valid_sync && !send_lreq_sync) || 
                             (csf_ctr == CSF_CYCLES-1) || 
                             send_ccomp || 
                             (send_lreq_sync && !lreq_sent && |stripe_valid);

      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          idle_frame_toggle <= #TCQ 1'b1;
        end else begin
          if (rand_df_reset)
            idle_frame_toggle <= #TCQ 1'b1;
          else if (rand_df_ctr == RAND_DF_MAX_CYCLES) 
            idle_frame_toggle <= #TCQ 1'b0;
        end
      end

      //Counter for the number of bytes in the rand data field of an idle
      //frame. This counter will reset at the start of an idle sequence after
      //valid data transmission, or whenever it reaches its max.  
      //The random data field can be between 509 and 515 bytes. 
      //Reset to 4 in the event a ccomp sequence started the idle and
      //therefore has 4 D0.0s inserted already. Plus two mask offs that may be
      //required
      //Reset to 2 in the event that only two mask offs are required 
      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          rand_df_ctr <= #TCQ 0;
        end else begin
          if (rand_df_reset)
            rand_df_ctr <= #TCQ (send_ccomp) ? (tx_idle2_selected ? IDLE2_CCOMP_CYCLES  : 
                                                                    IDLE1_CCOMP_CYCLES) : 2;
          else if (idle_frame_toggle)
            rand_df_ctr <= #TCQ rand_df_ctr + 1'b1;
        end
      end

      //*ASSERTION*
      // (ap_rand_df_ctr_overflows): The rand_df_ctr doesn't overflow

      //The Command and Status field counter.  This counter will start at
      //0 after the random data field is transmitted.  Otherwise the
      //idle_frame_toggle switch will indicate when it reaches CSF_CYCLES-1
      //and to stop counting.
      // Reset if:
      // 1. A clock compensation needs to be inserted
      // 2. Valid data is incoming
      wire reset_csf_ctr = send_ccomp || |stripe_valid || mask_idles;

      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          csf_ctr <= #TCQ CSF_CYCLES;
        end else begin
          if (reset_csf_ctr)
            csf_ctr <= #TCQ CSF_CYCLES;
          else if (rand_df_ctr == RAND_DF_MAX_CYCLES) 
            csf_ctr <= #TCQ 0;
          else if (!idle_frame_toggle)
            csf_ctr <= #TCQ csf_ctr + 1'b1;
        end
      end

      //*ASSERTION*
      // (ap_csf_ctr_maxed): the csf_ctr does not count past the max value
      
      //Select the correct random data charater, when an A or M is not
      //indicated a D0_0 is always sent.
      for (i2r_ii=0; i2r_ii < GT_BYTES; i2r_ii=i2r_ii+1) begin: i2_rand_gen
        always @(*) begin
          //Only sent D0_0s if the CFSM is about to be transmitted 
          if (rand_df_ctr == RAND_DF_MAX_CYCLES) begin 
            i2_rand[i2r_ii*8+:8]  = {GT_BYTES{D0_0}};
            i2_isk_rand[i2r_ii]   = {GT_BYTES{1'b0}};
          end else begin
            case ({i2_send_a[i2r_ii], i2_send_m[i2r_ii]})
              2'b10:  begin 
                i2_rand[i2r_ii*8+:8] = A_CHAR;
                i2_isk_rand[i2r_ii]  = 1'b1;
              end
              2'b01:  begin
                i2_rand[i2r_ii*8+:8] = M_CHAR;
                i2_isk_rand[i2r_ii]  = 1'b1;
              end
              default: begin 
                i2_rand[i2r_ii*8+:8] = D0_0;
                i2_isk_rand[i2r_ii]  = 1'b0;
              end
            endcase
          end
        end //end always
      end //end for (i2r_ii < GT_BYTES)

      //The Command and Status Field marker must be sent as the first 8 bytes
      //in the CS Field.  Two are sent per cycle.
      assign send_csfm = (csf_ctr < (8/GT_BYTES)) && !reset_csf_ctr;
      
      //Since the csf counter remains at a value of 20 when not in use we know
      //the CS Field needs to be transmitted whenever the value of the counter
      //is not 20
      assign send_csf  = (csf_ctr != CSF_CYCLES) && !reset_csf_ctr;
     
      //register the send_csf signal to be used in the scramblers to determine
      //if scrambling should be bypassed.
      //use the registered version in the scrambler since when send_csf
      //asserts it will pass through the lane_d stage before arriving to the
      //scrambler
      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          cs_field        <= #TCQ 0;
          cs_field_q      <= #TCQ 0;
          cs_field_start  <= #TCQ 0;
        end else begin 
          cs_field        <= #TCQ send_csf;
          cs_field_q      <= #TCQ (cs_field && !mask_idles);
          cs_field_start  <= #TCQ ((csf_ctr < (4/GT_BYTES)) && !mask_idles); // The M's
        end
      end

      //*COVERPOINT*
      // (cp_csf_terminated_after_csfm): a valid packet comes terminates the CSF directly 
      // after the cs field marker

      //*COVERPOINT*
      //(cp_csf_terminated_mid): the csf is terminated mid cs field

      //generate an idle for each lane
      for (i2_ii = 0; i2_ii < LINK_WIDTH; i2_ii=i2_ii+1) begin: idle2_lanes_gen
        //The appropriate data is selected for insertion into the idle stream.
        //This can be the clk comp seq, the cs field marker, the encoded cs
        //field, or the random data field.
        // Subtract two from the cs ctr to account for the csfm
        wire [7:0] csf_select                = tx_csf[i2_ii][(8-(csf_ctr-2)-1)*8+:8];
        assign     csf_select_encoded[i2_ii] = csencode(csf_select);

        //*ASSERTION*
        // (cp_csf_encoded_x): The csencode function must never result in X's

        always @(posedge gt_pcs_clk) begin
          if (gt_pcs_rst_q) begin
            idle2[i2_ii]     <= #TCQ 0;
            idle2_isk[i2_ii] <= #TCQ 0;
          end else begin
            if (send_ccomp) begin
              idle2[i2_ii]     <= #TCQ IDLE2_CCOMP_SEQ[(IDLE2_CCOMP_CYCLES-ccomp_ctr-1)*32+:32];
              idle2_isk[i2_ii] <= #TCQ IDLE2_CCOMP_SEQ_ISK[(IDLE2_CCOMP_CYCLES-ccomp_ctr-1)*4+:4];
            end else if (send_csfm) begin
              idle2[i2_ii]     <= #TCQ csfm[i2_ii][(CSM_CYCLES-csf_ctr-1)*GT_BYTES*8+:GT_BYTES*8];
              idle2_isk[i2_ii] <= #TCQ csfm_isk[(CSM_CYCLES-csf_ctr-1)*GT_BYTES+:GT_BYTES];
            end else if (send_csf) begin
              idle2[i2_ii]     <= #TCQ csf_select_encoded[i2_ii]; 
              idle2_isk[i2_ii] <= #TCQ 2'b00;
            end else begin
              idle2[i2_ii]     <= #TCQ i2_rand;
              idle2_isk[i2_ii] <= #TCQ i2_isk_rand;
            end
          end
        end
      end //end for (i2_ii < LINK_WIDTH)
    end //end if (IDLE2)
    else begin: no_idle2_seq_gen
      //Tie off these wires for the bind files
      assign i2_send_a = 0;
      assign i2_send_m = 0;
      assign send_csfm = 0;
      assign send_csf  = 0;
      assign send_ack  = 0;
      assign send_nack = 0;
      assign send_cmd  = 0;

      always @(posedge gt_pcs_clk) begin
        rand_df_ctr    <= #TCQ 0;
        i2_rand        <= #TCQ 0;
        i2_isk_rand    <= #TCQ 0;
        cs_field       <= #TCQ 0;
        cs_field_q     <= #TCQ 0;
        cs_field_start <= #TCQ 0;
      end
    end
  endgenerate
  // }}} IDLE2 Sequence Generator
  
  // {{{ IDLE Sequence Selector
  //Select the appropriate idle settings based on the parameters
  //or the tx_idle2_selected signal

  //*COVERPOINT*
  // (cp_idle2_selected): when both IDLE1 and IDLE2, the idle sequence selection logic pick both 
  // cases

  genvar sel_ii; //select 
  generate
    case ({(IDLE1 == 1), (IDLE2 == 1)})
      //IDLE1 Only mode
      {1'b1,1'b0}: begin: idle1_gen
        for (sel_ii = 0; sel_ii < LINK_WIDTH; sel_ii=sel_ii+1) begin: idle1_select_gen
          assign idle    [sel_ii] = idle1;
          assign idle_isk[sel_ii] = idle1_isk;
        end
      end

      //IDLE2 Only mode
      {1'b0,1'b1}: begin: idle2_gen
        for (sel_ii = 0; sel_ii < LINK_WIDTH; sel_ii=sel_ii+1) begin: idle2_select_gen
          assign idle    [sel_ii] = (mask_idles) ? {GT_BYTES{D0_0}} : idle2[sel_ii];
          assign idle_isk[sel_ii] = (mask_idles) ? {GT_BYTES{1'b0}} : idle2_isk[sel_ii];
        end 
      end

      //IDLE1 and IDLE 2 modes
      {1'b1,1'b1}: begin: idle1_idle2_gen
        for (sel_ii = 0; sel_ii < LINK_WIDTH; sel_ii=sel_ii+1) begin: idle1_idle2_select_gen
          assign idle    [sel_ii] = (tx_idle2_selected) ? 
                                    ((mask_idles) ? {GT_BYTES{D0_0}} : idle2[sel_ii]) : 
                                    idle1;
          assign idle_isk[sel_ii] = (tx_idle2_selected) ? 
                                    ((mask_idles) ? {GT_BYTES{1'b0}} : idle2_isk[sel_ii]) : 
                                    idle1_isk;
        end 
      end
    endcase
  endgenerate
  // }}} IDLE Sequence Selector
  
  // }}} + Idle Sequence Generator +------------

  // {{{ Sync Sequence Generator ------------
  //If IDLE2 mode is supported, generate the logic to create the
  //synchronization sequence.
  generate if (IDLE2) begin: sync_seq_gen
    //Define the synchronization sequence used in the descramblers
    //where the two LSB's is transmitted first
    reg   [2:0]             valid_cycles;
    reg   [GT_BYTES*8-1:0]  sync_seq_q;
    reg   [GT_BYTES-1:0]    sync_seq_isk_q;
    wire  [GT_BYTES-1:0]    sync_seq_isk_d;
    wire  [GT_BYTES*8-1:0]  sync_seq_d;
    wire                    drop_send_sync;
    wire  [2:0]             sync_seq_ctr_mod;

    //The Synchronization Sequence is (broken up by cycles): 
    //{MDDD, DMDD, DDMD, DDDM, DDDD}
    wire [159:0] SYNC_SEQ = {M_CHAR, D0_0,   D0_0,   D0_0,    // Cycle1
                             D0_0,   M_CHAR, D0_0,   D0_0,    // Cycle2
                             D0_0,   D0_0,   M_CHAR, D0_0,    // Cycle3
                             D0_0,   D0_0,   D0_0,   M_CHAR,  // Cycle4
                             D0_0,   D0_0,   D0_0,   D0_0};   // Cycle5

    //The sync seq isk wire marks the locations of the M_CHARs in the
    //SYNC_SEQ wire.
    wire [19:0] SYNC_SEQ_ISK = {4'b1000,  // Cycle1
                                4'b0100,  // Cycle2
                                4'b0010,  // Cycle3
                                4'b0001,  // Cycle4
                                4'b0000}; // Cycle5

    //Assert to send a link-request when a send_lreq_sync is available 
    //and the counter is less than the number of cycles it takes to
    //send the entrie sync squence.
    wire start_sync_sequence = (|tx_valid_sync && send_lreq_sync && (sync_seq_ctr < 4) && !lreq_sent && 
                                !indicate_lreq_sent) || 
                               (lreq_complete && early_lreq_sync);
    assign drop_send_sync = (sync_seq_ctr_mod == 4);

    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        send_sync <= #TCQ 0;
      end else begin
        if (drop_send_sync) begin
          send_sync <= #TCQ 0;
        end else if (start_sync_sequence) begin
          send_sync <= #TCQ 1;
        end
      end
    end

    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        valid_send_lreq <= #TCQ 0;
      end else begin
        if (lreq_complete && !early_lreq_sync) begin
          valid_send_lreq <= #TCQ 0;
        end else if (start_sync_sequence) begin
          valid_send_lreq <= #TCQ 1'b1;
        end
      end
    end

    //Count the number of cycles to transmit the synchronization
    //sequence and the valid data that follows.  This count should reset
    //when the link-request is done and increment as long as the
    //link-request is available indicated by sync_send
    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        sync_seq_ctr <= #TCQ 0;
      end else begin
        if (lreq_complete) begin
          sync_seq_ctr <= #TCQ 0;
        end else if (valid_send_lreq) begin
          sync_seq_ctr <= #TCQ sync_seq_ctr + 1'b1;
        end
      end
    end
      
    //*ASSERTION*
    //(ap_sync_seq_overflow): Sync sequence counter does not overflow

    //Based on the link width, the number of cycles to transmit the valid
    //link-request varies.  Done can not be asserted until all valid data
    //has been transmitted.
    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        valid_cycles <= #TCQ (LINK_WIDTH == 1) ? 2 : 
                             (LINK_WIDTH == 2) ? 1 : 
                                                 1;
      end else if (PPI_mode_1x) begin
        valid_cycles <= #TCQ 2;
      end else if (LINK_WIDTH == 2) begin
        valid_cycles <= #TCQ 1;
      end else if (LINK_WIDTH == 4) begin
        if (send_sync) begin
          valid_cycles <= #TCQ (shift_sync_seq) ? 0 : 1;
        end
      end
    end

    assign lreq_complete = (sync_seq_ctr == (SYNC_CYCLES-1)+valid_cycles);

    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        lreq_sent <= #TCQ 0;
      end else begin
        if (lreq_sent) begin
          lreq_sent <= #TCQ 1'b0;
        end else if (lreq_complete) begin
          lreq_sent <= #TCQ 1'b1;
        end
      end
    end

    //Indicate early to the ollm rx when the sync seq has been inserted 
    //to have new data by the time it actually completes. this is needed
    //since takes time to get synchronized
    assign indicate_lreq_complete = ((LINK_WIDTH == 1) || PPI_mode_1x) ? 
                                      (sync_seq_ctr == (SYNC_CYCLES-5)+valid_cycles) :
                                      (sync_seq_ctr == (SYNC_CYCLES-3)+valid_cycles);

    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        indicate_lreq_sent <= #TCQ 0;
      end else begin
        if (!send_lreq_sync) begin
          indicate_lreq_sent <= #TCQ 1'b0;
        end else if (indicate_lreq_complete || 
                    (lreq_complete && !indicate_lreq_sent && !early_lreq_sync)) begin
          indicate_lreq_sent <= #TCQ 1'b1;
        end
      end
    end
      
    // Register the send_lreq_sync signal for the lane_d logic to know when
    // to mask off the handshake data
    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        send_lreq_sync_q <= #TCQ 0;
      end else begin
        send_lreq_sync_q <= #TCQ send_lreq_sync;
      end
    end

    // For 4x modes, if there are two b2b LREQs to send, we may need to
    // shift the starting point of the SYNC since an LREQ only stripes
    // across 2 bytes and not the full 4 of the GT interface.
    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        shift_sync_seq <= #TCQ 0;
      end else if (!PPI_mode_1x && (LINK_WIDTH == 4) && !send_sync && lreq_complete) begin
        shift_sync_seq <= #TCQ (!shift_sync_seq) ? early_lreq_sync : 0;
      end 
    end

    // Wire the sync sequence to make selecting bytes/debug easier
    // Once it counts to the length of the sync sequence start back over at
    // 0. this is need for x4 cores with b2b lreqs
    assign sync_seq_ctr_mod = shift_sync_seq ? ((sync_seq_ctr+1)%5) : (sync_seq_ctr%5);
    assign sync_seq_d     = SYNC_SEQ[(SYNC_CYCLES-1-sync_seq_ctr_mod)*GT_BYTES*8+:GT_BYTES*8];
    assign sync_seq_isk_d = SYNC_SEQ_ISK[(SYNC_CYCLES-1-sync_seq_ctr_mod)*GT_BYTES+:GT_BYTES];

    assign sync_seq     = (shift_sync_seq) ? {sync_seq_q[15:0], sync_seq_d[31:16]}      : sync_seq_d;
    assign sync_seq_isk = (shift_sync_seq) ? {sync_seq_isk_q[1:0], sync_seq_isk_d[3:2]} : sync_seq_isk_d;

    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        sync_seq_q      <= #TCQ 0;
        sync_seq_isk_q  <= #TCQ 0;
      end else begin  
        sync_seq_q      <= #TCQ sync_seq_d;
        sync_seq_isk_q  <= #TCQ sync_seq_isk_d;
      end
    end

  end //end if (IDLE2)
  else begin: no_sync_seq_gen
    //Tie off signals not used in IDLE1 mode
    always @(posedge gt_pcs_clk) begin
      lreq_sent           <= #TCQ 0;
      indicate_lreq_sent  <= #TCQ 0;
      send_sync           <= #TCQ 0;
      send_lreq_sync_q    <= #TCQ 0;
      valid_send_lreq     <= #TCQ 0;
      shift_sync_seq      <= #TCQ 0;
      sync_seq_ctr        <= #TCQ 0;
    end
    assign sync_seq      = 0;
    assign sync_seq_isk  = 0;
    assign lreq_complete = 0;

  end endgenerate
  // }}} Sequence Selector Generator --------

  // {{{ Data Switch ------------------------
  //*ASSERTION*
  // (ap_lanes_equal): IDLE1/IDLE sequence is identical across all lanes
  // ignore lane comparison if there is valid data or the csfield
  genvar dsb_ii; // data switch bytes
  genvar dsl_ii; // data switch lanes

  //Select the correct data to output for each lane
  generate for (dsl_ii=0; dsl_ii < LINK_WIDTH; dsl_ii=dsl_ii+1) begin: data_switch_gen
    for (dsb_ii = 0; dsb_ii < GT_BYTES;  dsb_ii=dsb_ii+1) begin: ds_bytes_gen
      // No need to reset data bits
      always @(posedge gt_pcs_clk) begin
        //Always send the sync sequence first if there is one
        if (send_sync) begin
          lane_d  [dsl_ii][dsb_ii*8+:8] <= #TCQ sync_seq[dsb_ii*8+:8];
          lane_isk[dsl_ii][dsb_ii]      <= #TCQ sync_seq_isk[dsb_ii];
          lane_valid[dsl_ii][dsb_ii]    <= #TCQ 1'b1; 

        //Send any valid data
        end else begin
          // For a link width of 4 and IDLE2 mode, if a new LREQ needs to be sent right 
          // after the currently transmitting one we need to start the sync sequence on 
          // the lower two bytes after the last LREQ this is a special case required because 
          // if we are streaming LREQ/reset control symbols they must go out back to back
          if (lreq_complete && early_lreq_sync && (LINK_WIDTH == 4) && !PPI_mode_1x) begin
            // If an lreq just finished and another one if coming start the
            // SYNC sequence 
            if (!shift_sync_seq) begin
              lane_d  [dsl_ii][dsb_ii*8+:8] <= #TCQ (stripe_valid[dsb_ii]) ? stripe[dsl_ii][dsb_ii*8+:8] : 
                                                    (dsb_ii == 1)          ? M_CHAR :
                                                    (dsb_ii == 0)          ? D0_0   : 
                                                                             idle[dsl_ii][dsb_ii*8+:8];
              lane_isk[dsl_ii][dsb_ii]      <= #TCQ (stripe_valid[dsb_ii]) ? stripe_isk[dsl_ii][dsb_ii] :
                                                    (dsb_ii == 1)          ? 1'b1 :
                                                    (dsb_ii == 0)          ? 1'b0 : 
                                                                             idle_isk[dsl_ii][dsb_ii];
              lane_valid[dsl_ii][dsb_ii]    <= #TCQ 1'b1;
            end else begin
              lane_d  [dsl_ii][dsb_ii*8+:8] <= #TCQ (dsb_ii == 3)          ? D0_0 :
                                                    (dsb_ii == 2)          ? D0_0   : 
                                                    (stripe_valid[dsb_ii]) ? stripe[dsl_ii][dsb_ii*8+:8] :
                                                                             idle[dsl_ii][dsb_ii*8+:8];
              lane_isk[dsl_ii][dsb_ii]      <= #TCQ (dsb_ii == 3)          ? 1'b0 :
                                                    (dsb_ii == 2)          ? 1'b0   :
                                                    (stripe_valid[dsb_ii]) ? stripe_isk[dsl_ii][dsb_ii] :
                                                                             idle_isk[dsl_ii][dsb_ii];
              lane_valid[dsl_ii][dsb_ii]    <= #TCQ 1'b1;
            end
          end else begin
            lane_d  [dsl_ii][dsb_ii*8+:8] <= #TCQ (stripe_valid[dsb_ii]) ? stripe[dsl_ii][dsb_ii*8+:8] : 
                                                                           idle[dsl_ii][dsb_ii*8+:8];
            lane_isk[dsl_ii][dsb_ii]      <= #TCQ (stripe_valid[dsb_ii]) ? stripe_isk[dsl_ii][dsb_ii] :
                                                                           idle_isk[dsl_ii][dsb_ii];
            lane_valid[dsl_ii][dsb_ii]    <= #TCQ stripe_valid[dsb_ii];
          end
        end
      end //end always 
    end //end for (dsb_ii < GT_BYTES)
  end endgenerate

  //*COVERAGE*
  //(cp_lreq_b2b_in_4x):   Send out back to back lreqs in 4x mode
  //(cp_lreq_b2b_in_2x):   Send out back to back lreqs in 2x mode

  // }}} Data Switch ------------------------

  // {{{ Scramblers -------------------------
  //Generate a scrambler for each lane if the IDLE2 parameter is set

  //Declare those wires used only for the IDLE1 sequence generator.
  //These are created outside the scope of the generate in order to assist
  //in coverage in the bind files.  This enables automatic binding and
  //eliminates the need for heirarchical references.
  wire [GT_BYTES-1:0]   charisr       [LINK_WIDTH-1:0];
  wire [GT_BYTES-1:0]   bypass_scram  [LINK_WIDTH-1:0];

  genvar sb_ii;     // scrambler bypass
  genvar sxor_ii;   // scrambler xor 
  genvar sl_ii;     // scrambler lanes

  //If IDLE2 mode is supported then scramblers should be used for each lane
  generate if (IDLE2) begin: scrambler_gen
      for (sl_ii=0; sl_ii < LINK_WIDTH; sl_ii=sl_ii+1) begin: scram_lane_gen
        wire [(GT_BYTES*8)-1:0] scrambled_data;
        wire [16:0]             lfsr1_curr;
        wire [16:0]             lfsr2_curr;

        // *ASSERTION*
        // (ap_scrambler_charisr): In IDLE2 R's are only ever sent for the clk comp sequence
        // in which case data will always be aligned as charisr == 0111

        //Indicate if there is a K characer that is the special character R.
        //If so the LFSR must not be incremented
        assign charisr[sl_ii][0] = lane_isk[sl_ii][0] && (lane_d[sl_ii][7:0]   == R_CHAR);
        assign charisr[sl_ii][1] = lane_isk[sl_ii][1] && (lane_d[sl_ii][15:8]  == R_CHAR);
        assign charisr[sl_ii][2] = lane_isk[sl_ii][2] && (lane_d[sl_ii][23:16] == R_CHAR);
        assign charisr[sl_ii][3] = lane_isk[sl_ii][3] && (lane_d[sl_ii][31:24] == R_CHAR);

        wire [2:0] r_count = charisr[sl_ii][0] + charisr[sl_ii][1] + 
                             charisr[sl_ii][2] + charisr[sl_ii][3];

        // Scrambler to scrambler the first 16-bits in the 4 byte interface
        // This scrambler gets xor'd with the high bits of the data so we need
        // to pass it the high bits when looking for an R_CHAR
        srio_gen2_v4_1_16_oplm_lfsr #(
          .TCQ          (TCQ),
          .LANE         (sl_ii),    
          .SCRAMBLER    (1)
        ) oplm_lfsr1_tx_inst (   
          .gt_pcs_clk       (gt_pcs_clk),
          .gt_pcs_rst_q     (gt_pcs_rst_q),
          .load             (1'b0),
          .shift16_on_load  (1'b0),
          .load_value       (17'b0),
          .r_count          (r_count),  
          .lfsr_curr        (lfsr1_curr),
          .lfsr_8           () 
        );

        // Scrambler to scrambler the second 16-bits in the 4 byte interface
        // This scrambler gets xor'd with the low bits of the data so we need
        // to pass it the low bits when looking for an R_CHAR
        srio_gen2_v4_1_16_oplm_lfsr #(
          .TCQ          (TCQ),
          .LANE         (sl_ii),    
          .SCRAMBLER    (2)
        ) oplm_lfsr2_tx_inst (   
          .gt_pcs_clk       (gt_pcs_clk),
          .gt_pcs_rst_q     (gt_pcs_rst_q),
          .load             (1'b0),
          .shift16_on_load  (1'b0),
          .load_value       (17'b0),
          .r_count          (r_count),  
          .lfsr_curr        (lfsr2_curr),
          .lfsr_8           () 
        );

        //When scrambing the data the lfsr_scram uses a 1:17 methodology to
        //match the spec for bit "16" needs to be XORed with bit "15" of the
        //data since bit 15 will go out first.
        wire [31:0] lfsr_curr = {lfsr2_curr[15:0], lfsr1_curr[15:0]};

        for (sxor_ii = 0; sxor_ii < 32; sxor_ii=sxor_ii+1) begin: scrambled_data_xor_gen
          assign scrambled_data[31-sxor_ii] = lane_d[sl_ii][31-sxor_ii] ^ lfsr_curr[sxor_ii];
        end 
        
        //Check data bytes for scrambling. Scramble if:
        //1. not in the CS field
        //2. there is not valid data when scrambling is disabled through the cfg
        //3. there is not a k character
        //4. it is disabled by the parameter
        for (sb_ii=0; sb_ii < GT_BYTES; sb_ii=sb_ii+1) begin: bypass_scram_gen
          assign bypass_scram[sl_ii][sb_ii] = (cs_field_q && !lane_valid[sl_ii][sb_ii])       || 
                                              (PC_scram_disable && lane_valid[sl_ii][sb_ii])  ||
                                              lane_isk[sl_ii][sb_ii]                          || 
                                              (SCRAM == 0);
          //*COVERAGE*
          // (cp_bypass_scram): See all interesting combination of a scrambler bypass on 
          // idle sequences only

          //No need to have a reset on data bits
          always @(posedge gt_pcs_clk) begin
            //Pass on K characters
            scram_isk[sl_ii][sb_ii] <= #TCQ lane_isk[sl_ii][sb_ii];

            // Scrambler only non-K characters when idle2 is selected, otherwise passthrough
            if (bypass_scram[sl_ii][sb_ii] || !tx_idle2_selected_q) begin
              scram[sl_ii][sb_ii*8+:8] <= #TCQ lane_d[sl_ii][sb_ii*8+:8];
            end else begin 
              scram[sl_ii][sb_ii*8+:8] <= #TCQ scrambled_data[sb_ii*8+:8];
            end
          end //end always
        end //end for (sb_ii < GT_BYTES)
        
      end //end for (sl_ii < LANE_WIDTH)
    end //end if (IDLE2)
    else begin: no_scrambler_gen
      //Tie off these wires for the bind files
      for (sl_ii = 0; sl_ii < LINK_WIDTH; sl_ii=sl_ii+1) begin: noscram_lane_gen
        assign charisr[sl_ii]       = 0;
        assign bypass_scram[sl_ii]  = 0;

        always @* begin
          scram[sl_ii]     = lane_d[sl_ii];
          scram_isk[sl_ii] = lane_isk[sl_ii];
        end
      end //end for (sl_ii < LINK_WIDTH)
    end
  endgenerate
  // }}} Scramblers -------------------------

  // {{{ MGT Interface ----------------------
  // When in IDLE2 mode select the data output from the scramblers, otherwise
  // selected the data outputs from the data switch logic.
  genvar gtd_ii; // gt data _d
  generate for (gtd_ii=0; gtd_ii < LINK_WIDTH; gtd_ii=gtd_ii+1) begin: gttx_gen
    assign gttx_data_d[(gtd_ii*8*GT_BYTES)+:(8*GT_BYTES)] = scram[gtd_ii];
    assign gttx_charisk_d[(gtd_ii*GT_BYTES)+:GT_BYTES]    = scram_isk[gtd_ii];
  end endgenerate

  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      PPT_gttx_data    <= #TCQ 0;
      PPT_gttx_charisk <= #TCQ 0;
    end else begin
      PPT_gttx_data    <= #TCQ gttx_data_d;
      PPT_gttx_charisk <= #TCQ gttx_charisk_d;
    end
  end
  // }}} MGT Interface ----------------------

endmodule
// {{{ DISCLAIMER OF LIABILITY
//----------------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/phy/oplm/srio_gen2_v4_1_16_oplm_lfsr.v#3 $
//----------------------------------------------------------------------
//
// OPLM_LFSR
// Description:
// This module contains the logic to model an LFSR used in the 
// scrambler/descrambler of the OPLM.  This LFSR models the function
// f(x) = x^17 + x^8 + 1 
//
// Hierarchy:
// PHY_TOP
//    |___OPLM_TOP
//            |___OPLM_RX
//            |      |_____OPLM_LFSR <-- this module
//            |
//            |___OPLM_TX
//                   |_____OPLM_LFSR <-- this module
// ---------------------------------------------------------------------
`timescale 1ps/1ps

// ------------------------------------------------
// below attribute is added to supress the synthesis warnings in vivado tool 8:3332
(* DowngradeIPIdentifiedWarnings="yes" *)
// ------------------------------------------------

module srio_gen2_v4_1_16_oplm_lfsr #(
    parameter TCQ         = 100,
    parameter SHIFT_BITS  = 32,   // Shift by 16 or Shift by 32 bits.
    parameter LANE        = 0,    // Indicate which lane this is for the initial values
    parameter SCRAMBLER   = 0,    // Indicate if this is a scrambler, which one, 
                                  // or if 0 then its a descrambler
    parameter DESCRAMBLER = 0)    // Indicate if this is a descrambler, which one, 
                                  // or if 0 then its a descrambler                              
  (
    // {{{ port declarations ---------------
    // System Signals
    input               gt_pcs_clk,        //GT Clock
    input               gt_pcs_rst_q,      //GT reset
    input               load,              //load a new value into the LFSR
    input               shift16_on_load,   // Indicated if the load_value needs modification before loading
    input       [1:17]  load_value,        //new LFSR value
    input       [2:0]   r_count,           //Indicates number of 3's on this cycle
    output reg  [1:17]  lfsr_curr,         //LFSRs current value
    output reg  [1:17]  lfsr_8             //LFSRs current value shifted by 8
    // }}} end port declarations -----------
  );

  //Wire Declarations
  wire [1:17] shift_by_8;
  wire [1:17] shift_by_16;
  wire [1:17] shift_by_24;
  wire [1:17] shift_by_32;
  wire [1:17] load_value_mod;

  // {{{ Local Parameters
  // Local parameters for lfsr initialization taken from the PHY spec table 4-9
  // in the scrambling rules section 4.8.1.  Each value must have an offset of
  // 64 from any other init value.
  localparam LN0_INIT1 = 17'b1111_1111_1111_1111_1;
  localparam LN1_INIT1 = 17'b1111_1111_0000_0110_1;
  localparam LN2_INIT1 = 17'b0000_0000_1000_0110_1;
  localparam LN3_INIT1 = 17'b0000_0110_0111_1010_0;

  // If the scrambler is needed for the second 2 bytes in the 4 bytes gt interface
  // the init values need to start 16 shifts off from the first two bytes
  localparam LN0_INIT2 = 17'b1111_1111_0000_0000_1;
  localparam LN1_INIT2 = 17'b0000_1100_1111_0010_1;
  localparam LN2_INIT2 = 17'b0000_1100_0000_1101_0;
  localparam LN3_INIT2 = 17'b1111_1110_1111_0010_0;

  // Set the appropriate initial value based on the lane number
  // for the second scrambler/descrambler it needs to load the offset by 16-bit value
  localparam SCRAM_INIT = (LANE == 0 && (SCRAMBLER == 1 || DESCRAMBLER == 1)) ? LN0_INIT1 : 
                          (LANE == 1 && (SCRAMBLER == 1 || DESCRAMBLER == 1)) ? LN1_INIT1 :
                          (LANE == 2 && (SCRAMBLER == 1 || DESCRAMBLER == 1)) ? LN2_INIT1 :
                          (LANE == 3 && (SCRAMBLER == 1 || DESCRAMBLER == 1)) ? LN3_INIT1 :
                          (LANE == 0 && (SCRAMBLER == 2 || DESCRAMBLER == 2)) ? LN0_INIT2 : 
                          (LANE == 1 && (SCRAMBLER == 2 || DESCRAMBLER == 2)) ? LN1_INIT2 :
                          (LANE == 2 && (SCRAMBLER == 2 || DESCRAMBLER == 2)) ? LN2_INIT2 :
                          (LANE == 3 && (SCRAMBLER == 2 || DESCRAMBLER == 2)) ? LN3_INIT2 : 17'bX;
  // }}} end Local Parameters

  // {{{ shift_8(curr) function
  function [1:17] shift_8(
    input [1:17] curr_16,
    input [1:17] curr
  );
    begin
      shift_8 = {curr_16[9:16], curr[1:9]};
    end
  endfunction
  // }}} end shift_8

  // {{{ shift_16(curr) function
  // Calculate the next state for the LFSR when incrementing by 16-bits 
  // this increments as a parallelized form of the 17-bit polynomial 
  // f(x) = x^17 + x^8 + 1
  // Written as a function to be used multiple times with one code base.
  function [1:17] shift_16 (
    input [1:17] curr   //LFSR value to shift
  );
    begin
      shift_16[17] = curr[1];
      shift_16[16] = curr[17] ^ curr[8];
      shift_16[15] = curr[16] ^ curr[7];
      shift_16[14] = curr[15] ^ curr[6];
      shift_16[13] = curr[14] ^ curr[5];
      shift_16[12] = curr[13] ^ curr[4];
      shift_16[11] = curr[12] ^ curr[3];
      shift_16[10] = curr[11] ^ curr[2];
      shift_16[9]  = curr[10] ^ curr[1];
      shift_16[8]  = (curr[17] ^ curr[8]) ^ curr[9];
      shift_16[7]  = (curr[16] ^ curr[7]) ^ curr[8];
      shift_16[6]  = (curr[15] ^ curr[6]) ^ curr[7];
      shift_16[5]  = (curr[14] ^ curr[5]) ^ curr[6];
      shift_16[4]  = (curr[13] ^ curr[4]) ^ curr[5];
      shift_16[3]  = (curr[12] ^ curr[3]) ^ curr[4];
      shift_16[2]  = (curr[11] ^ curr[2]) ^ curr[3];
      shift_16[1]  = (curr[10] ^ curr[1]) ^ curr[2];
    end
  endfunction
  // }}} shift_16(curr) function

  // {{{ shift_24(curr) function
  // Calculate the next state for the LFSR when incrementing by 24-bits 
  // this increments as a parallelized form of the 17-bit polynomial 
  // f(x) = x^17 + x^8 + 1
  // Written as a function to be used multiple times with one code base.
  function [1:17] shift_24 (
    input [1:17] curr   //LFSR value to shift
  );
    begin
      shift_24[17] = curr[10] ^ curr[1];
      shift_24[16] = (curr[17] ^ curr[8]) ^ curr[9];
      shift_24[15] = (curr[16] ^ curr[7]) ^ curr[8];
      shift_24[14] = (curr[15] ^ curr[6]) ^ curr[7];
      shift_24[13] = (curr[14] ^ curr[5]) ^ curr[6];
      shift_24[12] = (curr[13] ^ curr[4]) ^ curr[5];
      shift_24[11] = (curr[12] ^ curr[3]) ^ curr[4];
      shift_24[10] = (curr[11] ^ curr[2]) ^ curr[3];
      shift_24[9]  = (curr[10] ^ curr[1]) ^ curr[2];
      shift_24[8]  = ((curr[17] ^ curr[8]) ^ curr[9]) ^ curr[1];  //17
      shift_24[7]  = ((curr[16] ^ curr[7]) ^ curr[8]) ^ (curr[17] ^ curr[8]); //18
      shift_24[6]  = ((curr[15] ^ curr[6]) ^ curr[7]) ^ (curr[16] ^ curr[7]); // 19
      shift_24[5]  = ((curr[14] ^ curr[5]) ^ curr[6]) ^ (curr[15] ^ curr[6]); // 20
      shift_24[4]  = ((curr[13] ^ curr[4]) ^ curr[5]) ^ (curr[14] ^ curr[5]); // 21
      shift_24[3]  = ((curr[12] ^ curr[3]) ^ curr[4]) ^ (curr[13] ^ curr[4]); // 22
      shift_24[2]  = ((curr[11] ^ curr[2]) ^ curr[3]) ^ (curr[12] ^ curr[3]); // 23
      shift_24[1]  = ((curr[10] ^ curr[1]) ^ curr[2]) ^ (curr[11] ^ curr[2]); // 24
    end
  endfunction
  // }}} shift_24(curr) function

  // {{{ shift_32(curr) function
  // Calculate the next state for the LFSR when incrementing by 32-bits 
  // this increments as a parallelized form of the 17-bit polynomial 
  // f(x) = x^17 + x^8 + 1
  // Written as a function to be used multiple times with one code base.
  function [1:17] shift_32 (
    input [1:17] curr   //LFSR value to shift
  );
    begin
      // Generate the function to shift by 32 bits (4 byte GT Interface)
      shift_32[17] = (curr[10] ^ curr[1]) ^ curr[2];
      shift_32[16] = ((curr[17] ^ curr[8]) ^ curr[9]) ^ curr[1];  //17
      shift_32[15] = ((curr[16] ^ curr[7]) ^ curr[8]) ^ (curr[17] ^ curr[8]); //18
      shift_32[14] = ((curr[15] ^ curr[6]) ^ curr[7]) ^ (curr[16] ^ curr[7]); // 19
      shift_32[13] = ((curr[14] ^ curr[5]) ^ curr[6]) ^ (curr[15] ^ curr[6]); // 20
      shift_32[12] = ((curr[13] ^ curr[4]) ^ curr[5]) ^ (curr[14] ^ curr[5]); // 21
      shift_32[11] = ((curr[12] ^ curr[3]) ^ curr[4]) ^ (curr[13] ^ curr[4]); // 22
      shift_32[10] = ((curr[11] ^ curr[2]) ^ curr[3]) ^ (curr[12] ^ curr[3]); // 23
      shift_32[9] = ((curr[10] ^ curr[1]) ^ curr[2]) ^ (curr[11] ^ curr[2]); // 24
      shift_32[8] = (((curr[17] ^ curr[8]) ^ curr[9]) ^ curr[1]) ^ (curr[10] ^ curr[1]); // 25
      shift_32[7] = (((curr[16] ^ curr[7]) ^ curr[8]) ^ (curr[17] ^ curr[8])) ^ ((curr[17] ^ curr[8]) ^ curr[9]); // 26
      shift_32[6] = (((curr[15] ^ curr[6]) ^ curr[7]) ^ (curr[16] ^ curr[7])) ^ ((curr[16] ^ curr[7]) ^ curr[8]); // 27
      shift_32[5] = (((curr[14] ^ curr[5]) ^ curr[6]) ^ (curr[15] ^ curr[6])) ^ ((curr[15] ^ curr[6]) ^ curr[7]); // 28
      shift_32[4] = (((curr[13] ^ curr[4]) ^ curr[5]) ^ (curr[14] ^ curr[5])) ^ ((curr[14] ^ curr[5]) ^ curr[6]); // 29
      shift_32[3] = (((curr[12] ^ curr[3]) ^ curr[4]) ^ (curr[13] ^ curr[4])) ^ ((curr[13] ^ curr[4]) ^ curr[5]); // 30
      shift_32[2] = (((curr[11] ^ curr[2]) ^ curr[3]) ^ (curr[12] ^ curr[3])) ^ ((curr[12] ^ curr[3]) ^ curr[4]); // 31
      shift_32[1] = (((curr[10] ^ curr[1]) ^ curr[2]) ^ (curr[11] ^ curr[2])) ^ ((curr[11] ^ curr[2]) ^ curr[3]); // 32
    end
  endfunction
  // }}} shift_32(curr) function

  // Calculate what an 8-bit shift would be since if a K character is present we need to skip it
  assign shift_by_8  = shift_8(shift_16(lfsr_curr), lfsr_curr);
  assign shift_by_16 = shift_16(lfsr_curr);
  assign shift_by_24 = shift_24(lfsr_curr);
  assign shift_by_32 = shift_32(lfsr_curr);

  // If we are loading new data we need to check if there should be a 16-bit shift on the load
  // value before it is loaded. This will occur if an M is detected such that the two bytes
  // to load were from a previous cycle and so the load_value requires more than just a 32 bit shift
  // to get back in sync with the data.
  assign load_value_mod = shift16_on_load ? shift_16(load_value) : load_value;

  //Do not increment the LFSR for R characters.
  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      lfsr_curr <= #TCQ SCRAM_INIT;

    end else begin
      //For descramblers enable loading a new value into the LFSR
      if (((DESCRAMBLER == 1) || (DESCRAMBLER == 2)) && load) begin
        // Shift it once to be in line with the next incoming data
        // to remain in sync with the incoming data, the load value must be shifted by one cycle
        // If this is descrambler 2, then it needs to be offset by 16 bits from lfsr 1
        lfsr_curr <= #TCQ (DESCRAMBLER == 1) ? shift_32(load_value_mod) : 
                          (DESCRAMBLER == 2) ? shift_32(shift_16(load_value_mod)) : 17'bX;

      end else begin
        //If there is an R figure out how much to shift by
        case (r_count)
          // Full Shift (32)
          0: begin
            lfsr_curr <= #TCQ shift_by_32;
            lfsr_8    <= #TCQ shift_8(shift_16(shift_by_32), shift_by_32);
          end
          // Shift by 24
          1: begin
            lfsr_curr <= #TCQ shift_by_24;
            lfsr_8    <= #TCQ shift_8(shift_16(shift_by_24), shift_by_24);
          end
          // Shift by 16
          2: begin
            lfsr_curr <= #TCQ shift_by_16;
            lfsr_8    <= #TCQ shift_8(shift_16(shift_by_16), shift_by_16);
          end
          // Shift by 8
          3: begin
            lfsr_curr <= #TCQ shift_by_8;
            lfsr_8    <= #TCQ shift_8(shift_16(shift_by_8), shift_by_8);
          end
          // No Shift
          4: begin
            lfsr_curr <= #TCQ lfsr_curr;
            lfsr_8    <= #TCQ lfsr_8;
          end
          // Invalid R count
          default: begin
            lfsr_curr <= #TCQ 17'bX;
            lfsr_8    <= #TCQ 17'bX;
          end
        endcase
      end
    end
  end

endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/phy/oplm/srio_gen2_v4_1_16_oplm_top.v#1 $
//----------------------------------------------------------------------
//
// OPLM_TOP
// Description:
// This module instantiates all the submodules of the OPLM design
//
// Hierarchy:
// PHY_TOP
//    |___OPLM_TOP <-- this module
//
// ---------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_oplm_top
  #(
    parameter TCQ           = 100,
    parameter LINK_WIDTH    = 1,                     // {1, 2, 4}
    parameter GT_BYTES      = 4,                     // GT Interface Bytes
    parameter DEBUG         = 0,                     // GT Interface Bytes
    parameter DATA_WIDTH    = LINK_WIDTH*GT_BYTES*8, // Data width
    parameter CHARIS_WIDTH  = LINK_WIDTH*GT_BYTES,   // Charisk bus width
    parameter IDLE1         = 1,                     // {0, 1}
    parameter IDLE2         = 0,                     // {0, 1}
    parameter MODE_XG       = 5,                     // {1, 2, 3, 5, 6}
    parameter SCRAM         = 0,                     // {0, 1}
    parameter GT_REG        = 1,                     // {0, 1} Register GT inputs
    parameter SIM_TRAIN     = 0,                     // {0: FULL, 1: DIVIDED TIMERS}     
    parameter EVAL          = 1)                     // Evaluation Core
  (
    // {{{ port declarations ---------------
    // System Signals
    input                             gt_pcs_clk,             //GT Clock /2
    input                             gt_pcs_rst,             //GT Clock /2 Reset
    input                             phy_clk,                //PHY Clock
    input                             phy_rst,                //PHY Clock Reset
    input                             sim_train_en,           //Enables the sim_train parameter

    // User Global Signals
    input                             UG_force_reinit,        //Forces link only rst

    // OLLM TX Interface
    input   [63:0]                    PT_tx_data,             //Transmit Data
    input   [7:0]                     PT_tx_charisk,          //Character is K
    input   [1:0]                     PT_tx_valid,            //Valid
    input                             PT_tx_early_lreq,       //One cycle early LREQ indicator
    input                             PT_ccomp_grant,         //Clock Comp. Granted
    input                             PT_send_lreq,           //Link Request

    output reg                        PP_port_initialized,    //Port Initialized
    output                            PP_ccomp_req,           //Clock Comp. Request
    output reg                        PP_idle2_selected,      //IDLE2 Sequence Sel.
    output reg                        PP_idle_selected,       //IDLE Sequence Sel.
    output                            PP_lreq_sent,           //Link Request Done

    // OLLM RX Interface
    output  [63:0]                    PP_rx_data,             //Receive Data
    output  [7:0]                     PP_rx_charisk,          //Character is K
    output  [1:0]                     PP_rx_valid,            //Valid
    output                            PP_out_of_sync,         //Descram Out of Sync
    output reg                        PP_mode_1x = 0,         //In 1x mode

    // MGT TX Interface
    output  [DATA_WIDTH-1:0]          PP_gttx_data,           //Transmit Data 
    output  [CHARIS_WIDTH-1:0]        PP_gttx_charisk,        //Character is K
    output  [LINK_WIDTH-1:0]          PP_gttx_inhibit,        //TX inhibit

    // MGT RX Interface
    input   [DATA_WIDTH-1:0]          GT_gtrx_data,           //Receive Data
    input   [CHARIS_WIDTH-1:0]        GT_gtrx_charisk,        //Character is K
    input   [CHARIS_WIDTH-1:0]        GT_gtrx_chariscomma,    //Character is Comma
    input   [CHARIS_WIDTH-1:0]        GT_gtrx_disperr,        //Disperity Error
    input   [CHARIS_WIDTH-1:0]        GT_gtrx_notintable,     //Not in Table
    input   [LINK_WIDTH-1:0]          GT_gtrx_chanisaligned,  //Channel is Aligned
    input                             GT_gtrx_reset_req,      //RX Buffer Error
    input   [LINK_WIDTH-1:0]          GT_gtrx_reset_done,     //Resets are done.
    output                            PP_gtrx_reset,          //Reset the RX Buffers
    output                            PP_gtrx_chanbonden,     //Enable Chanel Bonding
    output reg                        PP_rx_lane_r,           //LaneR is the Master

    // PHY Config Interface
    input                             PC_scram_disable,       //Scrambler Disable
    input   [2:0]                     PC_force_lane,          //Force train down
    input                             PC_port_disable,        //Disable link init.
    input                             PC_idle2_enable,        //Enable IDLE2 mode forced

    output  [LINK_WIDTH-1:0]          PP_rx_scram_en,         //scram enabled on rx
    output  [LINK_WIDTH-1:0]          PP_receiver_trained,    //trained indicator
    output  [LINK_WIDTH-1:0]          PP_idle2_rcvd,          //CS field of the IDLE2 Sequence detected
    output  [LINK_WIDTH*4-1:0]        PP_rx_lane_number,      //RX lane number 
    output  [LINK_WIDTH*3-1:0]        PP_rx_port_width,       //RX active port width 
    output  [LINK_WIDTH*GT_BYTES-1:0] PP_gt_decode_error,     //GT error detected 
    output  [LINK_WIDTH-1:0]          PP_lane_sync,           //lane sync status

    // PHY Equalization Interface
    input   [LINK_WIDTH-1:0]          PE_gttx_cmd,            // Command to send in the CSF
    input   [LINK_WIDTH*2-1:0]        PE_gttx_tap_m1_cmd,     // Tap -1 Command
    input   [LINK_WIDTH*2-1:0]        PE_gttx_tap_p1_cmd,     // Tap +1 Command
    input   [LINK_WIDTH-1:0]          PE_gttx_reset_emphasis, // Cmd Reset Emphasis
    input   [LINK_WIDTH-1:0]          PE_gttx_preset_emphasis,// Cmd Preset Emphasis
    input   [LINK_WIDTH*2-1:0]        PE_gttx_tap_m1_status,  // Current Tap -1 Status
    input   [LINK_WIDTH*2-1:0]        PE_gttx_tap_p1_status,  // Current Tap +1 Status
    input   [LINK_WIDTH-1:0]          PE_gttx_ack,            // Recieved cmd was ACK'd
    input   [LINK_WIDTH-1:0]          PE_gttx_nack,           // Recieved cmd was NACK'd

    output   [LINK_WIDTH-1:0]         PP_gtrx_cmd,            // Command recieved in the CSF
    output   [LINK_WIDTH*2-1:0]       PP_gtrx_tap_m1_cmd,     // Tap -1 Command
    output   [LINK_WIDTH*2-1:0]       PP_gtrx_tap_p1_cmd,     // Tap +1 Command
    output   [LINK_WIDTH-1:0]         PP_gtrx_reset_emphasis, // Cmd Reset Emphasis
    output   [LINK_WIDTH-1:0]         PP_gtrx_preset_emphasis,// Cmd Preset Emphasis
    output   [LINK_WIDTH*2-1:0]       PP_gtrx_tap_m1_status,  // Current Tap -1 Status of link partner
    output   [LINK_WIDTH*2-1:0]       PP_gtrx_tap_p1_status,  // Current Tap +1 Status of link partner
    output   [LINK_WIDTH-1:0]         PP_gtrx_ack,            // Sent cmd was ACK'd
    output   [LINK_WIDTH-1:0]         PP_gtrx_nack,           // Sent cmd was NACK'd

    output  [95:0]                    PP_debug                //Debug Port with cfg register values
    // }}} end port declarations -----------
  );

// added below macro to fix the CR# 735137
// synthesis translate_off 
  // {{{ Catch Bad Parameters
  //Catch any invalid parameter conditions
  initial begin
    if ((LINK_WIDTH == 3) || (LINK_WIDTH > 5)) begin
      $display("ERROR: Invalid Link Width Setting. LINK_WIDTH=%0d", LINK_WIDTH);
      $finish;
    end
    if (!IDLE2 && (MODE_XG > 5)) begin
      $display("ERROR: Invalid Combination of IDLE modes and Speed. IDLE2=%0d MODE_XG=%0d", 
               IDLE2, MODE_XG);
      $finish;
    end
    if (!IDLE1 && (MODE_XG <= 5)) begin
      $display("ERROR: Invalid Combination of IDLE modes and Speed. IDLE1=%0d MODE_XG=%0d", 
               IDLE1, MODE_XG);
      $finish;
    end
    if (IDLE1 && (MODE_XG == 6)) begin
      $display("ERROR: Cannot use IDLE1 mode in a 6G configuration.");
      $finish;
    end
    if ((MODE_XG == 4) || (MODE_XG > 6)) begin
      $display("ERROR: Invalid Speed Setting. MODE_XG=%0d", MODE_XG);
      $finish;
    end
  end
  // }}}
// synthesis translate_on

  // {{{ Wire Declarations -----------------
  wire                      PPI_port_initialized;    
  wire                      PPR_idle2_selected;    
  wire                      PPR_idle_selected;    
  wire                      PPI_mode_1x;

  //Registered GT RX Signals for the OPLM RX
  wire [DATA_WIDTH-1:0]     PPG_gtrx_data;         
  wire [CHARIS_WIDTH-1:0]   PPG_gtrx_chariskchar;      
  wire [CHARIS_WIDTH-1:0]   PPG_gtrx_charisa;      
  wire [CHARIS_WIDTH-1:0]   PPG_gtrx_charisk;      
  wire [CHARIS_WIDTH-1:0]   PPG_gtrx_charisr;      
  wire [CHARIS_WIDTH-1:0]   PPG_gtrx_charism;      
  wire [CHARIS_WIDTH-1:0]   PPG_gtrx_charispd;      
  wire [CHARIS_WIDTH-1:0]   PPG_gtrx_charissc;      
  wire [CHARIS_WIDTH-1:0]   PPG_gtrx_chariscomma;  
  wire [CHARIS_WIDTH-1:0]   PPG_gtrx_invalid;      
  wire [LINK_WIDTH-1:0]     PPG_gtrx_chanisaligned;
  wire                      PPG_gtrx_reset_req;    
  wire [LINK_WIDTH-1:0]     PPG_gtrx_reset_done;   

  //Additional Debug Signals
  wire                      PPI_n_lanes_aligned;   
  wire                      PPI_n_lanes_rdy;       
  wire                      PPI_x1_mode_detected;  
  wire [3:0]                PPI_init_state;
  wire                      PPI_reinit_sm;
  wire                      PPI_idle_select_en;
  wire                      PPI_rx_lane_r;

  // Debug Bus assignment
  // The debug bus provides as output to chipscope those signals that may be 
  // useful for debugging link bring up. 
  // These are not registered output because of this.
  assign PP_debug[0]      = PPR_idle2_selected;
  assign PP_debug[1]      = PP_mode_1x;
  assign PP_debug[2]      = PPR_idle_selected;
  assign PP_debug[3]      = PPI_port_initialized;
  assign PP_debug[4]      = PP_rx_lane_r;
  assign PP_debug[5]      = PP_gtrx_chanbonden;
  assign PP_debug[9:6]    = 4'b0;
  assign PP_debug[13:10]  = PPG_gtrx_chanisaligned;
  assign PP_debug[29:14]  = PPG_gtrx_chariscomma;
  assign PP_debug[33:30]  = PP_gttx_inhibit;
  assign PP_debug[34]     = PPG_gtrx_reset_req;
  assign PP_debug[35]     = PPI_n_lanes_aligned;
  assign PP_debug[36]     = PPI_n_lanes_rdy;
  assign PP_debug[37]     = PPI_x1_mode_detected;
  assign PP_debug[41:38]  = PPI_init_state;
  assign PP_debug[42]     = PP_out_of_sync;
  assign PP_debug[48:43]  = 0;
  // }}} Wire Declarations -----------------

  // {{{ Register Reset for Fanout ---------
  reg gt_pcs_rst_q = 1;
  reg phy_rst_q     = 1;

  always @(posedge gt_pcs_clk) begin
    gt_pcs_rst_q <= #TCQ gt_pcs_rst;
  end

  always @(posedge phy_clk) begin
    phy_rst_q <= #TCQ phy_rst;
  end
  // }}}------------------------------------

  // {{{ oplm_gtregisters inst
  //--------------------------------------------
  srio_gen2_v4_1_16_oplm_gtregisters
    #(.TCQ                       (TCQ),
      .LINK_WIDTH                (LINK_WIDTH),
      .GT_BYTES                  (GT_BYTES),
      .GT_REG                    (GT_REG))
    oplm_gtregisters_inst
     (.gt_pcs_clk                (gt_pcs_clk),
      .gt_pcs_rst_q              (gt_pcs_rst_q),
      .GT_gtrx_data              (GT_gtrx_data),
      .GT_gtrx_charisk           (GT_gtrx_charisk),
      .GT_gtrx_chariscomma       (GT_gtrx_chariscomma),
      .GT_gtrx_disperr           (GT_gtrx_disperr),
      .GT_gtrx_notintable        (GT_gtrx_notintable),
      .GT_gtrx_chanisaligned     (GT_gtrx_chanisaligned),
      .GT_gtrx_reset_req         (GT_gtrx_reset_req),
      .GT_gtrx_reset_done        (GT_gtrx_reset_done),
      .PPG_gtrx_data             (PPG_gtrx_data),
      .PPG_gtrx_chariskchar      (PPG_gtrx_chariskchar),
      .PPG_gtrx_charisa          (PPG_gtrx_charisa),
      .PPG_gtrx_charisk          (PPG_gtrx_charisk),
      .PPG_gtrx_charisr          (PPG_gtrx_charisr),
      .PPG_gtrx_charism          (PPG_gtrx_charism),
      .PPG_gtrx_charispd         (PPG_gtrx_charispd),
      .PPG_gtrx_charissc         (PPG_gtrx_charissc),
      .PPG_gtrx_chariscomma      (PPG_gtrx_chariscomma),
      .PPG_gtrx_invalid          (PPG_gtrx_invalid),
      .PPG_gtrx_chanisaligned    (PPG_gtrx_chanisaligned),
      .PPG_gtrx_reset_req        (PPG_gtrx_reset_req),
      .PPG_gtrx_reset_done       (PPG_gtrx_reset_done));
  // }}} End oplm_gtregisters inst

  // {{{ oplm_tx inst ----------------------
  // Instantiate the TX path for the OPLM
  srio_gen2_v4_1_16_oplm_tx
  #(
    .TCQ         (TCQ),
    .LINK_WIDTH  (LINK_WIDTH),
    .GT_BYTES    (GT_BYTES),
    .IDLE1       (IDLE1),
    .IDLE2       (IDLE2),
    .MODE_XG     (MODE_XG),
    .SCRAM       (SCRAM),
    .EVAL        (EVAL)
  ) oplm_tx_inst (
    .gt_pcs_clk              (gt_pcs_clk),
    .gt_pcs_rst_q            (gt_pcs_rst_q),
    .phy_clk                 (phy_clk),
    .phy_rst_q               (phy_rst_q),
    .PT_tx_data              (PT_tx_data),
    .PT_tx_charisk           (PT_tx_charisk),
    .PT_tx_valid             (PT_tx_valid),
    .PT_tx_early_lreq        (PT_tx_early_lreq),
    .PT_ccomp_grant          (PT_ccomp_grant),
    .PT_send_lreq            (PT_send_lreq),
    .PPT_ccomp_req           (PP_ccomp_req),
    .PPT_lreq_sent           (PP_lreq_sent),
    .PPT_gttx_data           (PP_gttx_data),
    .PPT_gttx_charisk        (PP_gttx_charisk),
    .PE_gttx_cmd             (PE_gttx_cmd), 
    .PE_gttx_tap_m1_cmd      (PE_gttx_tap_m1_cmd),
    .PE_gttx_tap_p1_cmd      (PE_gttx_tap_p1_cmd),
    .PE_gttx_reset_emphasis  (PE_gttx_reset_emphasis),
    .PE_gttx_preset_emphasis (PE_gttx_preset_emphasis),
    .PE_gttx_tap_m1_status   (PE_gttx_tap_m1_status),
    .PE_gttx_tap_p1_status   (PE_gttx_tap_p1_status),
    .PE_gttx_ack             (PE_gttx_ack),
    .PE_gttx_nack            (PE_gttx_nack), 
    .PC_scram_disable        (PC_scram_disable),
    .PPI_port_initialized    (PPI_port_initialized),
    .PPR_idle_selected       (PPR_idle_selected),
    .PPR_idle2_selected      (PPR_idle2_selected),
    .PPI_mode_1x             (PPI_mode_1x),
    .PPI_lane_sync           (PP_lane_sync));
  // }}} -----------------------------------

  // {{{ oplm_init inst --------------------
  // Instantiate port initialization state machines
  srio_gen2_v4_1_16_oplm_init 
  #(
    .TCQ           (TCQ),
    .MODE_XG       (MODE_XG),
    .LINK_WIDTH    (LINK_WIDTH),
    .GT_BYTES      (GT_BYTES),
    .IDLE1         (IDLE1),
    .IDLE2         (IDLE2),
    .SIM_TRAIN     (SIM_TRAIN)
  ) oplm_init_inst (
    .gt_pcs_clk            (gt_pcs_clk),
    .gt_pcs_rst_q          (gt_pcs_rst_q),
    .sim_train_en           (sim_train_en),
    .UG_force_reinit        (UG_force_reinit),
    .PC_force_lane          (PC_force_lane),
    .PC_port_disable        (PC_port_disable),
    .PPR_idle_selected      (PPR_idle_selected),
    .PPG_gtrx_charispd      (PPG_gtrx_charispd),
    .PPG_gtrx_charissc      (PPG_gtrx_charissc),
    .PPG_gtrx_charisa       (PPG_gtrx_charisa),
    .PPG_gtrx_chariscomma   (PPG_gtrx_chariscomma),
    .PPG_gtrx_invalid       (PPG_gtrx_invalid),
    .PPG_gtrx_chanisaligned (PPG_gtrx_chanisaligned),
    .PPG_gtrx_reset_req     (PPG_gtrx_reset_req),
    .PPG_gtrx_reset_done    (PPG_gtrx_reset_done),
    .PPI_mode_1x            (PPI_mode_1x),
    .PPI_rx_lane_r          (PPI_rx_lane_r),
    .PPI_lane_sync          (PP_lane_sync),
    .PPI_port_initialized   (PPI_port_initialized),
    .PPI_reinit_sm          (PPI_reinit_sm),
    .PPI_idle_select_en     (PPI_idle_select_en),
    .PPI_gtrx_reset         (PP_gtrx_reset),
    .PPI_gtrx_chanbonden    (PP_gtrx_chanbonden),
    .PPI_gttx_inhibit       (PP_gttx_inhibit),
    .PPI_n_lanes_aligned    (PPI_n_lanes_aligned),
    .PPI_n_lanes_rdy        (PPI_n_lanes_rdy),
    .PPI_x1_mode_detected   (PPI_x1_mode_detected),
    .PPI_init_state         (PPI_init_state));  
  // }}} -----------------------------------
    
  // {{{ oplm_rx inst ----------------------
  // Instantiate the RX path of the OPLM
  srio_gen2_v4_1_16_oplm_rx
  #(
    .TCQ        (TCQ),
    .LINK_WIDTH (LINK_WIDTH),
    .GT_BYTES   (GT_BYTES),
    .DEBUG      (DEBUG),
    .IDLE1      (IDLE1),
    .IDLE2      (IDLE2),
    .MODE_XG    (MODE_XG),
    .SCRAM      (SCRAM)
   ) oplm_rx_inst (
    .gt_pcs_clk              (gt_pcs_clk),              
    .gt_pcs_rst_q            (gt_pcs_rst_q),
    .phy_clk                  (phy_clk),
    .phy_rst_q                (phy_rst_q),
    .PPR_rx_data              (PP_rx_data),
    .PPR_rx_charisk           (PP_rx_charisk),
    .PPR_rx_valid             (PP_rx_valid),
    .PPR_out_of_sync          (PP_out_of_sync),
    .PPG_gtrx_data            (PPG_gtrx_data),
    .PPG_gtrx_chariskchar     (PPG_gtrx_chariskchar),
    .PPG_gtrx_charisk         (PPG_gtrx_charisk),
    .PPG_gtrx_charisr         (PPG_gtrx_charisr),
    .PPG_gtrx_charism         (PPG_gtrx_charism),
    .PPG_gtrx_charispd        (PPG_gtrx_charispd),
    .PPG_gtrx_charissc        (PPG_gtrx_charissc),
    .PPG_gtrx_invalid         (PPG_gtrx_invalid),
    .PC_scram_disable         (PC_scram_disable), 
    .PPR_receiver_trained     (PP_receiver_trained),    
    .PPR_rx_lane_number       (PP_rx_lane_number),    
    .PPR_rx_port_width        (PP_rx_port_width),    
    .PPR_rx_scram_en          (PP_rx_scram_en),
    .PPR_gt_decode_error      (PP_gt_decode_error),
    .PPR_idle2_rcvd           (PP_idle2_rcvd),
    .PPR_gtrx_cmd             (PP_gtrx_cmd), 
    .PPR_gtrx_tap_m1_cmd      (PP_gtrx_tap_m1_cmd),
    .PPR_gtrx_tap_p1_cmd      (PP_gtrx_tap_p1_cmd),
    .PPR_gtrx_reset_emphasis  (PP_gtrx_reset_emphasis),
    .PPR_gtrx_preset_emphasis (PP_gtrx_preset_emphasis),
    .PPR_gtrx_tap_m1_status   (PP_gtrx_tap_m1_status),
    .PPR_gtrx_tap_p1_status   (PP_gtrx_tap_p1_status),
    .PPR_gtrx_ack             (PP_gtrx_ack),
    .PPR_gtrx_nack            (PP_gtrx_nack),
    .PPI_port_initialized     (PPI_port_initialized),
    .PPI_reinit_sm            (PPI_reinit_sm),
    .PPI_idle_select_en       (PPI_idle_select_en),
    .PPI_mode_1x              (PPI_mode_1x),
    .PPI_rx_lane_r            (PPI_rx_lane_r),
    .PPI_lane_sync            (PP_lane_sync),
    .PC_idle2_enable          (PC_idle2_enable),
    .PPR_idle_selected        (PPR_idle_selected),
    .PPR_idle2_selected       (PPR_idle2_selected));
  // }}} -----------------------------------

  // {{{ Sync outputs that are also shared in the oplm
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin 
      PP_idle2_selected   <= #TCQ IDLE2;
      PP_idle_selected    <= #TCQ (IDLE2 ^ IDLE1);
      PP_mode_1x          <= #TCQ (LINK_WIDTH == 1);
      PP_port_initialized <= #TCQ 0;
      PP_rx_lane_r        <= #TCQ 0;
    end else begin
      PP_idle2_selected   <= #TCQ PPR_idle2_selected;
      PP_idle_selected    <= #TCQ PPR_idle_selected;
      PP_mode_1x          <= #TCQ PPI_mode_1x;
      PP_port_initialized <= #TCQ PPI_port_initialized;
      PP_rx_lane_r        <= #TCQ PPI_rx_lane_r;
    end
  end
  // }}} end sync

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/phy/oplm/srio_gen2_v4_1_16_eval_gt_pcs_clk.v#1 $
//----------------------------------------------------------------------
//
// EVAL_GT_PCS_CLK
// Description:
// This is the evaluation timer for the PHY TX which runs on the gt_pcs_clk
//
// Hierarchy:
// PHY_TOP
//    |___OPLM_TOP
//            |___OPLM_TX
//                    |___EVAL_GT_PCS_CLK <-- this module
// ---------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_eval_gt_pcs_clk #(
  parameter TCQ     = 100,
  parameter MODE_XG = 5)  // Line rates {1/1.25, 2/2.5, 3/3.125, 5/5, 6/6.25}
(
  output reg  flag  = 0,
  input       rst,
  input       clk
);

  //This clock will operate in the GT_PCS_CLK domain. Based on the selected mode,
  //the timeout will be calculated to obtain a time of 8 hours.
  //MODE_XG | GT_PCS_CLK (Mhz)  | Period (us) | Cycle Count Needed      
  //   1    |    31.25          |  .032       |   900,000,000,000,000 ~ (255^6)*3  = 7.3 hrs
  //   2    |    62.5           |  .016       | 1,800,000,000,000,000 ~ (255^6)*7  = 8.5 hrs
  //   3    |    78.13          |  .0123      | 2,341,463,414,634,146 ~ (255^6)*9  = 8.4 hrs
  //   5    |    125            |  .008       | 3,600,000,000,000,000 ~ (255^6)*13 = 7.9 hrs
  //   6    |    156.25         |  .0064      | 4,500,000,000,000,000 ~ (255^6)*16 = 7.8 hrs

  // Need 5 Stages reguardless of mode (A-E)
  // Initialize all registers to 0 since no reset is attached to this module

  // Stage A
  //------------------------------
  reg   [7:0] a = 0;
  reg         a_out = 0;
  wire        a_ceo;
  wire        a_en;

  assign a_en = 1'b1;

  always @(posedge clk) begin 
    if (rst) begin
      a     <= #TCQ 0;
      a_out <= #TCQ 0;
    end else begin
      if (a_en) begin
        a   <= #TCQ a + 1;
      end
      a_out <= #TCQ a_ceo;
    end
  end

  assign a_ceo = a_en & (&a);

  // Stage B
  //------------------------------
  reg   [7:0] b = 0;
  reg         b_out = 0;
  wire        b_ceo;
  wire        b_en;

  assign b_en = a_out;

  always @(posedge clk) begin
    if (rst) begin
      b     <= #TCQ 0;
      b_out <= #TCQ 0;
    end else begin
      if (b_en) begin
        b   <= #TCQ b + 1;
      end
      b_out <= #TCQ b_ceo;
    end
  end

  assign b_ceo = b_en & (&b);


  // Stage C
  //------------------------------
  reg   [7:0] c = 0;
  reg         c_out = 0;
  wire        c_ceo;
  wire        c_en;

  assign c_en = b_out;

  always @(posedge clk) begin
    if (rst) begin
      c     <= #TCQ 0;
      c_out <= #TCQ 0;
    end else begin
      if (c_en) begin
        c   <= #TCQ c + 1;
      end
      c_out <= #TCQ c_ceo;
    end
  end

  assign c_ceo = c_en & (&c);


  // Stage D
  //------------------------------
  reg   [7:0] d = 0;
  reg         d_out = 0;
  wire        d_ceo;
  wire        d_en;

  assign d_en = c_out;

  always @(posedge clk) begin
    if (rst) begin
      d     <= #TCQ 0;
      d_out <= #TCQ 0;
    end else begin
      if (d_en) begin
        d   <= #TCQ d + 1;
      end
      d_out <= #TCQ d_ceo;
    end
  end

  assign d_ceo = d_en & (&d);


  // Stage E
  //------------------------------
  reg   [7:0] e = 0;
  reg         e_out = 0;
  wire        e_ceo;
  wire        e_en;

  assign e_en = d_out;

  always @(posedge clk) begin
    if (rst) begin
      e     <= #TCQ 0;
      e_out <= #TCQ 0;
    end else begin
      if (e_en) begin
        e   <= #TCQ e + 1;
      end
      e_out <= #TCQ e_ceo;
    end
  end

  assign e_ceo = e_en & (&e);

  // Stage F
  // -----------------------------
  //This clock will operate in the GT_PCS_CLK domain. Based on the selected mode,
  //the timeout will be calculated to obtain a time of 8 hours.
  //MODE_XG | GT_PCS_CLK (Mhz)  | Period (us) | Cycle Count Needed      
  //   1    |    31.25          |  .032       |   900,000,000,000,000 ~ (255^6)*3  = 7.3 hrs
  //   2    |    62.5           |  .016       | 1,800,000,000,000,000 ~ (255^6)*7  = 8.5 hrs
  //   3    |    78.13          |  .0123      | 2,341,463,414,634,146 ~ (255^6)*9  = 8.4 hrs
  //   5    |    125            |  .008       | 3,600,000,000,000,000 ~ (255^6)*13 = 7.9 hrs
  //   6    |    156.25         |  .0064      | 4,500,000,000,000,000 ~ (255^6)*16 = 7.8 hrs
 
  //Figure out the number to count to on the last stage based on the mode
  //calculations
  localparam LAST_STAGE_COUNT = (MODE_XG == 1) ? 3 :
                                (MODE_XG == 2) ? 7 :
                                (MODE_XG == 3) ? 9 :
                                (MODE_XG == 5) ? 13 : 16;
  reg  [4:0]  f = 0;
  wire        f_ceo;
  wire        f_en;

  assign f_en = e_out;

  always @(posedge clk) begin
    if (rst) begin
      f <= #TCQ 0;
    end else begin
      if (f_en) begin
        f <= #TCQ f + 1;
      end
    end
  end

  assign f_ceo = f_en & (f == LAST_STAGE_COUNT);

  // Generate the expire flag
  //------------------------------
  always @(posedge clk) begin
    if (rst) begin
      flag <= #TCQ 0;

    end else if (f_ceo) begin
      flag <= #TCQ 1;
    end
  end

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/phy/oplm/srio_gen2_v4_1_16_oplm_rx.v#4 $
//----------------------------------------------------------------------
//
// OPLM_RX
// Description:
// This module is the RX path of the OPLM.  It is responsible for the
// following:
// 1. Receiving Data from the link partner from the GTs
// 2. Descrambling Data if IDLE2 mode is selected
// 3. Destriping the data if the link width is > 1 indication it was striped
// 4. Aligning data as necessary.
// 5. Decoding the IDLE2 sequence is selected and providing the necessary
//    Data to the configuration registers
//
// Hierarchy:
// PHY_TOP
//    |___OPLM_TOP
//            |___OPLM_RX <-- this module
// --------------------------------------------------------------------
`timescale 1ps/1ps

// ------------------------------------------------
// below attribute is added to supress the synthesis warnings in vivado tool 8:3332
(* DowngradeIPIdentifiedWarnings="yes" *)
// ------------------------------------------------

module srio_gen2_v4_1_16_oplm_rx
  #(
    parameter TCQ           = 100,
    parameter LINK_WIDTH    = 1,                     // {1, 2, 4}
    parameter GT_BYTES      = 4,                     // Bytes on the GT interface per lane
    parameter DEBUG         = 0,                     // Bytes on the GT interface per lane
    parameter DATA_WIDTH    = LINK_WIDTH*GT_BYTES*8, // Incoming Data width
    parameter CHARIS_WIDTH  = LINK_WIDTH*GT_BYTES,   // Incoming Charisk bus width
    parameter IDLE1         = 1,                     // {0, 1}
    parameter IDLE2         = 0,                     // {0, 1}
    parameter MODE_XG       = 5,                     // {1, 2, 3, 5, 6}
    parameter SCRAM         = 0)                     // {0, 1}
  (
    // {{{ port declarations ---------------
    // System Signals
    input                                 gt_pcs_clk,             //GT Clock
    input                                 gt_pcs_rst_q,           //GT Clock Reset
    input                                 phy_clk,                 //Phy Clock 
    input                                 phy_rst_q,               //Phy Reset 

    // OPLM Synchronization Interface
    output reg  [63:0]                    PPR_rx_data,             //Aligned data
    output reg  [7:0]                     PPR_rx_charisk,          //Aligned data
    output reg  [1:0]                     PPR_rx_valid,            //Valid
    output reg                            PPR_out_of_sync,         //Descrams out of sync

    // MGT RX Interface
    input       [DATA_WIDTH-1:0]          PPG_gtrx_data,           //Receive Data
    input       [CHARIS_WIDTH-1:0]        PPG_gtrx_chariskchar,    //Character is K
    input       [CHARIS_WIDTH-1:0]        PPG_gtrx_charisk,        //Character is /K/
    input       [CHARIS_WIDTH-1:0]        PPG_gtrx_charisr,        //Character is /R/
    input       [CHARIS_WIDTH-1:0]        PPG_gtrx_charism,        //Character is /M/
    input       [CHARIS_WIDTH-1:0]        PPG_gtrx_charispd,       //Character is /PD/
    input       [CHARIS_WIDTH-1:0]        PPG_gtrx_charissc,       //Character is /SC/
    input       [CHARIS_WIDTH-1:0]        PPG_gtrx_invalid,        //Disperity Error/Not in Table
    
    // PHY Config Interface
    input                                 PC_scram_disable,        //Scrambler Disable
    output reg  [LINK_WIDTH-1:0]          PPR_receiver_trained,    //Received Trained
    output reg  [LINK_WIDTH*4-1:0]        PPR_rx_lane_number,      //RX lanes number
    output reg  [LINK_WIDTH*3-1:0]        PPR_rx_port_width,       //RX active port width
    output reg  [LINK_WIDTH-1:0]          PPR_rx_scram_en,         //Receivers Scram EN
    output reg  [LINK_WIDTH*GT_BYTES-1:0] PPR_gt_decode_error,     //8B/10B GT Error
    output reg  [LINK_WIDTH-1:0]          PPR_idle2_rcvd,          //the idle2 CSFM was recieved
   
    // PHY Equalization Interface
    output reg  [LINK_WIDTH-1:0]          PPR_gtrx_cmd,            // Command recieved in the CSF
    output reg  [LINK_WIDTH*2-1:0]        PPR_gtrx_tap_m1_cmd,     // Tap -1 Command
    output reg  [LINK_WIDTH*2-1:0]        PPR_gtrx_tap_p1_cmd,     // Tap +1 Command
    output reg  [LINK_WIDTH-1:0]          PPR_gtrx_reset_emphasis, // Cmd Reset Emphasis
    output reg  [LINK_WIDTH-1:0]          PPR_gtrx_preset_emphasis,// Cmd Preset Emphasis
    output reg  [LINK_WIDTH*2-1:0]        PPR_gtrx_tap_m1_status,  // Current Tap -1 Status of link partner
    output reg  [LINK_WIDTH*2-1:0]        PPR_gtrx_tap_p1_status,  // Current Tap +1 Status of link partner
    output reg  [LINK_WIDTH-1:0]          PPR_gtrx_ack,            // Sent cmd was ACK'd
    output reg  [LINK_WIDTH-1:0]          PPR_gtrx_nack,           // Sent cmd was NACK'd

    //OPLM Internal Signals
    input                                 PPI_port_initialized,    //link is init.
    input                                 PPI_reinit_sm,           //Re-initialize
    input                                 PPI_idle_select_en,      //Look for the idle seq 
    input                                      PPI_mode_1x,             //Mode 1x Selected
    input                                      PPI_rx_lane_r,           //1x on lane R
    input       [LINK_WIDTH     -1:0]          PPI_lane_sync,           //Lanes Sync'd
    input                                      PC_idle2_enable,         //Force IDLE2
    output reg                                 PPR_idle_selected,       //idle seq selected
    output reg                                 PPR_idle2_selected       //idle2 selected
    // }}} end port declara     tions -----------
  );

  // {{{ Wire Declarations      -----------------

  wire  [(GT_BYTES*8)-1:0]       rx_data_exp           [LINK_WIDTH-1:0];
  reg   [(GT_BYTES*8)-1:0]       rx_data_exp_q         [LINK_WIDTH-1:0];
  wire  [GT_BYTES-1:0]           rx_chariskchar_exp    [LINK_WIDTH-1:0];
  reg   [GT_BYTES-1:0]           rx_chariskchar_exp_q  [LINK_WIDTH-1:0];
  wire  [GT_BYTES-1:0]           rx_charisk_exp        [LINK_WIDTH-1:0];
  wire  [GT_BYTES-1:0]           rx_charisr_exp        [LINK_WIDTH-1:0];
  wire  [GT_BYTES-1:0]           rx_charism_exp        [LINK_WIDTH-1:0];
  wire  [GT_BYTES-1:0]           rx_charispdsc_exp     [LINK_WIDTH-1:0];
  wire  [GT_BYTES-1:0]           rx_invalid_exp        [LINK_WIDTH-1:0];

  // Descrambling 
  reg   [(GT_BYTES*8)-1:0]       descram            [LINK_WIDTH-1:0];
  reg   [GT_BYTES-1:0]           descram_isk        [LINK_WIDTH-1:0];
  reg   [GT_BYTES-1:0]           descram_invalid    [LINK_WIDTH-1:0];
  reg   [GT_BYTES-1:0]           descram_pd_sc      [LINK_WIDTH-1:0];
  reg   [LINK_WIDTH-1:0]         ln_out_of_sync;
  reg                       gt_out_of_sync;

  // CS Field
  wire  [GT_BYTES-1:0]      cs_field;
  reg   [3:0]               cs_ctr;
  reg                       cs_ctr_en;
  reg                       cs_ctr_en_q;
  reg                       cs_ctr_en_qq;
  reg                       cs_ctr_en_qqq;
  wire  [GT_BYTES-1:0]      cs_start_d;
  reg   [GT_BYTES-1:0]      cs_start;
  reg   [GT_BYTES-1:0]      cs_start_q;
  reg                       cs_aligned_q;
  wire  [GT_BYTES-1:0]      cs_interrupt;

  //Destriping Logic Signals
  wire  [DATA_WIDTH-1:0]    destripe_gen;
  wire  [CHARIS_WIDTH-1:0]  destripe_isk_gen;
  wire  [CHARIS_WIDTH-1:0]  destripe_invalid_gen;
  wire  [CHARIS_WIDTH-1:0]  destripe_pdsc_gen;

  reg   [DATA_WIDTH-1:0]    destripe_q;
  reg   [CHARIS_WIDTH-1:0]  destripe_isk_q;
  reg   [CHARIS_WIDTH-1:0]  destripe_invalid_q;
  reg   [3:0]               destripe_pdsc_q; // originally CHARIS_WIDTH, reduced to remove warning

  //Byte alignment Signals
  reg   [3:0]               byte_alignment;
  reg   [3:0]               byte_alignment_q;
  reg   [1:0]               aligned_start_idx_1x;
  reg   [1:0]               aligned_end_idx_1x;
  reg   [2:0]               aligned_start_idx_2x;
  reg   [2:0]               aligned_end_idx_2x;
  wire  [2:0]               aligned_start_idx_2x_lower;
  wire  [2:0]               aligned_end_idx_2x_lower;
  wire                      csymbol_start_2x;
  wire                      csymbol_end_2x;
  reg                       csymbol_monitor;
  reg                       csymbol_toggle_q;
  reg                       csymbol_toggle_qq;
  wire                      correct_byte_alignment_1x;
  wire                      correct_byte_alignment;
  wire                      multiple_alignments;
  reg   [3:0]               upper_byte_alignment;
  wire  [3:0]               realign;
  wire                      valid_realign;
  reg                       flush_stored_q;
  reg                       realign_allowed_q;
  reg                       new_byte_alignment_q;
  reg   [3:0]               locked_bytes;
  reg   [9:0]               byte1_stored;
  reg   [9:0]               byte2_stored;
  reg   [9:0]               byte3_stored;


  // Shared across x4 and x2 modes
  reg [63:0]                gt_rx_data_nx_q;
  reg [7:0]                 gt_rx_charisk_nx_q;
  reg [1:0]                 gt_rx_valid_nx_q;
  
  // Only for a x4 trained core
  reg [63:0]                gt_rx_data_q;
  reg [7:0]                 gt_rx_charisk_q;
  reg [3:0]                 gt_rx_valid_q;

  reg [63:0]                gt_rx_data_1x_q;
  reg [7:0]                 gt_rx_charisk_1x_q;
  reg [1:0]                 gt_rx_valid_1x_q;

  reg  [10:0]      byte_alignment_2x_d;
  reg              csymbol_monitor_2x;
  reg  [6:0]      byte_alignment_1x_d;



  reg   [DATA_WIDTH-1:0]    destripe;
  
  reg   [CHARIS_WIDTH-1:0]  destripe_isk;

  reg   [CHARIS_WIDTH-1:0]  destripe_invalid;
  
  reg   [CHARIS_WIDTH-1:0]  destripe_pdsc;
  // Clock Domain Crossing signals
  reg [DATA_WIDTH-1:0]      gt_rx_data;
  reg [CHARIS_WIDTH-1:0]    gt_rx_charisk;
  reg [CHARIS_WIDTH-1:0]    gt_rx_valid;
  reg [2:0]      rx_1x_align_next_state;
  reg [2:0]      rx_1x_align_state;
  reg  [2:0]      rx_align_next_state;
  
  reg  [2:0]      rx_align_state;


  generate if (DEBUG == 1)
    begin: extra_debug_signals_on
         (* mark_debug = "true" *)
         wire   [DATA_WIDTH-1:0]    debug_destripe = destripe;
         
         (* mark_debug = "true" *)
         wire   [CHARIS_WIDTH-1:0]  debug_destripe_isk = destripe_isk;

         (* mark_debug = "true" *)
         wire   [CHARIS_WIDTH-1:0]  debug_destripe_invalid = destripe_invalid;
         
         (* mark_debug = "true" *)
         wire   [CHARIS_WIDTH-1:0]  debug_destripe_pdsc = destripe_pdsc;
         // Clock Domain Crossing signals
         (* mark_debug = "true" *)
         wire [DATA_WIDTH-1:0]      debug_gt_rx_data = gt_rx_data;
         (* mark_debug = "true" *)
         wire [CHARIS_WIDTH-1:0]    debug_gt_rx_charisk = gt_rx_charisk;
         (* mark_debug = "true" *)
         wire [CHARIS_WIDTH-1:0]    debug_gt_rx_valid = gt_rx_valid;
         (* mark_debug = "true" *)
         wire [2:0]      debug_rx_1x_align_next_state = rx_1x_align_next_state;
         (* mark_debug = "true" *)
         wire [2:0]      debug_rx_1x_align_state = rx_1x_align_state;
         (* mark_debug = "true" *)
         wire  [2:0]      debug_rx_align_next_state = rx_align_next_state;
         
         (* mark_debug = "true" *)
         wire  [2:0]      debug_rx_align_state = rx_align_state;
    end
  endgenerate



//RX 1X State Machine States
  localparam ALIGN_1X           = 10'd0;
  localparam ONE_BIT_SHIFT      = 10'd1;
  localparam TWO_BIT_SHIFT      = 10'd2;
  localparam THREE_BIT_SHIFT    = 10'd3;
  localparam INTER_STATE        = 10'd4;
  localparam INTER_STATE2       = 10'd5;
  localparam INTER_STATE1       = 10'd6;
  
//RX 1X logic signals
  reg csymbol_monitor_1x;
  reg upper_nibble_pd;
  reg lower_nibble_pd;
  reg upper_nibble_pd_q;
  reg lower_nibble_pd_q;
  reg fresh_pd;
  reg stale_pd;
  

  reg start_1x_transaction;

  // }}} Wire Declarations -----------------

  // {{{ Local Parameters ------------------

  // SRIO Protocol Parameters
  // -------------------------
  // The redundancy lane
  localparam R = (LINK_WIDTH == 2) ? 1 : 
                 (LINK_WIDTH == 4) ? 2 : 0; 
  
  //Parameters for the CS Field Marker Encodings (table 4-8 of PHY spec)
  localparam DECODE_00 = 8'h67;  //D7.3 character
  localparam DECODE_01 = 8'h78;  //D24.3 character
  localparam DECODE_10 = 8'h7E;  //D30.3 character
  localparam DECODE_11 = 8'hF8;  //D24.7 character

  // Need an inverted decode as well for the CS field
  localparam INV_DECODE_11 = 8'h98;  //~D7.3 character
  localparam INV_DECODE_10 = 8'h87;  //~D24.3 character
  localparam INV_DECODE_01 = 8'h81;  //~D30.3 character
  localparam INV_DECODE_00 = 8'h07;  //~D24.7 character


  //Start of packet K characters used for alignment
  localparam PD_CHAR = 8'h7C;
  localparam SC_CHAR = 8'h1C;

  // Inserted characters for realignment
  localparam R_CHAR  = 8'hFD;
  localparam D0_0    = 8'h00;

  //OPLM RX Defined Parameters
  //--------------------------
  //The length of the CS Field minus the MMMM markers in cycles
  // 32-bits *2 for check bits = 64-bits
  // 64-bits encoded as 2 bits eq 1 byte, 64/2= 32 bytes
  // 32 bytes + 4 for the second half of the marker == 40 bytes
  localparam CS_BYTES  = 40;
  localparam CS_CYCLES = CS_BYTES/GT_BYTES; // 10 cyles;

  //The number of possible lanes
  localparam VALID_LANES = 4;

  // }}} Local Parameters ------------------

  // {{{ MGT Interface ---------------------
  //Expand the gtrx_data bus out into a two dimensional array to easily
  //access throughout this module
  genvar exp_ii; // expand 
  generate
    for (exp_ii=0; exp_ii < LINK_WIDTH; exp_ii=exp_ii+1) begin: expand_rx_data_gen
      assign rx_data_exp[exp_ii]        = PPG_gtrx_data[(exp_ii*GT_BYTES*8)+:(GT_BYTES*8)];
      assign rx_chariskchar_exp[exp_ii] = PPG_gtrx_chariskchar[(exp_ii*GT_BYTES)+:GT_BYTES];
      assign rx_charisk_exp[exp_ii]     = PPG_gtrx_charisk[(exp_ii*GT_BYTES)+:GT_BYTES];
      assign rx_charisr_exp[exp_ii]     = PPG_gtrx_charisr[(exp_ii*GT_BYTES)+:GT_BYTES];
      assign rx_charism_exp[exp_ii]     = PPG_gtrx_charism[(exp_ii*GT_BYTES)+:GT_BYTES];
      assign rx_charispdsc_exp[exp_ii]  = PPG_gtrx_charispd[(exp_ii*GT_BYTES)+:GT_BYTES] | 
                                          PPG_gtrx_charissc[(exp_ii*GT_BYTES)+:GT_BYTES];
      assign rx_invalid_exp[exp_ii]     = PPG_gtrx_invalid[(exp_ii*GT_BYTES)+:GT_BYTES];

      // Pass on any GT errors to the PHY Cfg space
      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          PPR_gt_decode_error[(exp_ii*GT_BYTES)+:GT_BYTES] <= #TCQ 0;

        // Only start monitoring for errors after the port is initialized
        end else if (!PPI_port_initialized) begin
          PPR_gt_decode_error[(exp_ii*GT_BYTES)+:GT_BYTES] <= #TCQ 0;
        
        end else begin
          PPR_gt_decode_error[(exp_ii*GT_BYTES)+:GT_BYTES] <= #TCQ rx_invalid_exp[exp_ii];
        end
      end //end always
    end // end for (exp_ii < LINK_WIDTH)
  endgenerate
  // }}} MGT Interface ---------------------

  // {{{ Idle Sequence Detector ------------
  //Declare those wires used only for the IDLE1 sequence detector.
  //These are created outside the scope of the generate in order to assist
  //in coverage in the bind files.  This enables automatic binding and
  //eliminates the need for heirarchical references.
  wire sync_lost;
  wire sync_lost_ln0;
  wire sync_lost_ln_r;

  //When both idle modes are supported, generate the sequence detection logic.
  generate
    if (IDLE1 && IDLE2) begin: idle_seq_select_gen
      reg  [2:0]              charisk_ctr;
      reg  [1:0]              charisd_ctr;
      wire                    sync_aquired;
      reg                     sync_aquired_q;
      reg  [LINK_WIDTH-1:0]   lane_sync_q;

      //Register lane_sync to be used to check for when sync switches lanes
      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          lane_sync_q <= #TCQ 0;
        end else begin
          lane_sync_q <= #TCQ PPI_lane_sync;
        end
      end

      //Monitor lane 0 and lane R for lane synchronization. Once sync is 
      //obtained that lane can be monitored for the idle sequence
      assign sync_lost_ln0  = (lane_sync_q[0] & ~PPI_lane_sync[0]);
      assign sync_lost_ln_r = (lane_sync_q[R] & ~PPI_lane_sync[R]);

      //*COVERAGE*
      //(cp_sync_lost_0): Sync is lost on lane 0

      //*COVERAGE*
      //(cp_sync_lost_r): Sync is lost on lane R

      assign sync_aquired   = PPI_lane_sync[0] | PPI_lane_sync[R];
      assign sync_lost      = (sync_aquired_q & ~sync_aquired) | sync_lost_ln0 | sync_lost_ln_r;

      //*COVERPOINT*
      //(cp_sync_switch_0): Lane sync is on lane 0 then switches to lane R to triggeer a sync lost

      //*ASSERTION*
      //(ap_sync_switch_detected_0): when a lane sync switches from lane 0 to R a switch is 
      //detected and sync is lost.

      //*COVERPOINT*
      //(cp_sync_switch_r): Lane sync is on lane R then switches to lane 0 to triggeer a sync lost
      
      //*ASSERTION*
      //(ap_sync_switch_detected_r): when a lane sync switches from lane 0 to R a switch is
      //detected and sync is lost.
      
      //*COVERPOINT*
      //(cp_sync_lost): Lane sync is aquired then lost before idle is selected

      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          sync_aquired_q <= #TCQ 1'b0;
        end else begin 
          sync_aquired_q <= #TCQ sync_aquired;
        end
      end

      //When sync is aquired monitor the lane for K charateres.  When 16
      //K characters are detected consecutively, IDLE1 mode is used.
      //Alignment should not matter at this point, so we will just count
      //two K characters at a time and reset if two are not seen
      wire idle_select_enable = sync_aquired && !PPR_idle_selected && PPI_idle_select_en;

      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          charisk_ctr <= #TCQ 0;
        end else begin 
          if (sync_lost || PPI_reinit_sm) begin
            charisk_ctr <= #TCQ 0;

          //count the number of K character received on the monitored lane
          end else if (idle_select_enable) begin
            //Monitoriing on lane 0
            if (PPI_lane_sync[0]) begin
              if (&rx_chariskchar_exp[0]) begin
                charisk_ctr <= #TCQ charisk_ctr + 1'b1;
              end else begin
                charisk_ctr <= #TCQ 0;
              end

            //Monitoring on lane R
            end else begin
              if (&rx_chariskchar_exp[R]) begin
                charisk_ctr <= #TCQ charisk_ctr + 1'b1;
              end else begin
                charisk_ctr <= #TCQ 0;
              end
            end
          end
        end
      end

      //When sync is aquired monitor the lane for D charateres.  When 8
      //D characters are detected consecutively, IDLE2 mode is used.
      //Alignment should not matter at this point, 8 should be seen in either
      //case
      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          charisd_ctr <= #TCQ 0;
        end else begin 
          if (sync_lost || PPI_reinit_sm) begin
            charisd_ctr <= #TCQ 0;

          //count the number of D character received on the monitored lane
          end else if (idle_select_enable) begin
            //Monitoring on lane 0
            if (PPI_lane_sync[0]) begin
              if (!(&rx_chariskchar_exp[0])) begin
                charisd_ctr <= #TCQ charisd_ctr + 1'b1;
              end else begin
                charisd_ctr <= #TCQ 0;
              end

            //Monitoring on lane R
            end else begin
              if (!(&rx_chariskchar_exp[R])) begin
                charisd_ctr <= #TCQ charisd_ctr + 1'b1;
              end else begin
                charisd_ctr <= #TCQ 0;
              end
            end
          end
        end
      end

      //*COVERPOINT*/
      //(cp_idle2_selected):IDLE1 and IDLE2 come up with both idle1 selected and idle2 selected

      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          PPR_idle_selected   <= #TCQ 0;
          PPR_idle2_selected  <= #TCQ IDLE2;
        end else begin
          // If the initialization state machines need to start over, reset
          // these ports
          if (PPI_reinit_sm) begin
            PPR_idle_selected   <= #TCQ 0;
            PPR_idle2_selected  <= #TCQ IDLE2;

          // If the CSRs disabled IDLE2 selection, ignore the counters
          end else if (!PC_idle2_enable && !PPI_port_initialized && PPI_idle_select_en) begin
            PPR_idle_selected   <= #TCQ 1'b1;
            PPR_idle2_selected  <= #TCQ 1'b0;
           
          // Look for 4 cycles of k-chars's for ILDE1 mode,
          // Look for 2 cycles of D0.0's for IDLE2 mode
          end else if (charisk_ctr[2] || charisd_ctr[1]) begin
            PPR_idle_selected   <= #TCQ 1'b1;
            PPR_idle2_selected  <= #TCQ charisd_ctr[1];
          end
        end
      end
    end else if (IDLE1) begin: idle1_only_select_gen
      //For IDLE1 only mode, tie off the idle being selected
      always @(posedge gt_pcs_clk) begin
        PPR_idle_selected  <= #TCQ 1'b1; 
        PPR_idle2_selected <= #TCQ 1'b0;
      end
      
      //Tie off these signals for bind files
      assign sync_lost      = 0;
      assign sync_lost_ln0  = 0;
      assign sync_lost_ln_r = 0;
    
    end else if (IDLE2) begin: idle2_only_select_gen
      //For IDLE2 only mode, tie off the idle being selected
      always @(posedge gt_pcs_clk) begin
        PPR_idle_selected  <= #TCQ 1'b1; 
        PPR_idle2_selected <= #TCQ 1'b1; 
      end

      //Tie off these signals for bind files
      assign sync_lost      = 0;
      assign sync_lost_ln0  = 0;
      assign sync_lost_ln_r = 0;
    end //end if (IDLE2)
  endgenerate
  // }}} Idle Sequence Detector ------------

  // {{{ Command and Status Decoder --------
  // For IDLE2 mode, generate the detection logic to decode the commmand and
  // status field of the idle sequence.  For IDLE1 this field does not exist
  genvar cs_ii;
  generate
    if (IDLE2) begin: cs_decoder_gen
      // {{{ CSDECODE Function
      //the csdeencode function deencodes the CS Field using 16 bits at a time 
      //to create a 2-bit value as indicated by the PHY Spec in table 4-8
      function [7:0] csdecode (
        input [31:0] x //value to decode
      );
        begin
          case(x[7:0])
            DECODE_00, INV_DECODE_00: csdecode[1:0] = 2'b00;
            DECODE_01, INV_DECODE_01: csdecode[1:0] = 2'b01;
            DECODE_10, INV_DECODE_10: csdecode[1:0] = 2'b10;
            DECODE_11, INV_DECODE_11: csdecode[1:0] = 2'b11;
            default:   csdecode[1:0] = 2'bXX;
          endcase
          case(x[15:8])
            DECODE_00, INV_DECODE_00: csdecode[3:2] = 2'b00;
            DECODE_01, INV_DECODE_01: csdecode[3:2] = 2'b01;
            DECODE_10, INV_DECODE_10: csdecode[3:2] = 2'b10;
            DECODE_11, INV_DECODE_11: csdecode[3:2] = 2'b11;
            default:   csdecode[3:2] = 2'bXX;
          endcase
          case(x[23:16])
            DECODE_00, INV_DECODE_00: csdecode[5:4] = 2'b00;
            DECODE_01, INV_DECODE_01: csdecode[5:4] = 2'b01;
            DECODE_10, INV_DECODE_10: csdecode[5:4] = 2'b10;
            DECODE_11, INV_DECODE_11: csdecode[5:4] = 2'b11;
            default:   csdecode[5:4] = 2'bXX;
          endcase
          case(x[31:24])
            DECODE_00, INV_DECODE_00: csdecode[7:6] = 2'b00;
            DECODE_01, INV_DECODE_01: csdecode[7:6] = 2'b01;
            DECODE_10, INV_DECODE_10: csdecode[7:6] = 2'b10;
            DECODE_11, INV_DECODE_11: csdecode[7:6] = 2'b11;
            default:   csdecode[7:6] = 2'bXX;
          endcase
        end
      endfunction
      // }}} CSDECODE Function
      
      // For each lane sample the CS Field 
      for (cs_ii = 0; cs_ii < LINK_WIDTH; cs_ii = cs_ii+1) begin: cs_ln_decode
        wire [7:0] decode_1000; // various alignments of the cs field decoded
        wire [7:0] decode_0100;
        wire [7:0] decode_0010;
        wire [7:0] decode_0001;

        reg        sample_csf_data;
        reg [63:0] rx_csf;
        reg [2:0]  rx_port_width;
        reg [3:0]  rx_lane_number;

        // decode the cs field for when in arrives on a two byte alignment or
        // shifted by one byte.
        assign decode_1000 = csdecode(rx_data_exp[cs_ii]);
        assign decode_0100 = csdecode({rx_data_exp_q[cs_ii][23:0],rx_data_exp[cs_ii][31:24]});
        assign decode_0010 = csdecode({rx_data_exp_q[cs_ii][15:0],rx_data_exp[cs_ii][31:16]});
        assign decode_0001 = csdecode({rx_data_exp_q[cs_ii][7:0],rx_data_exp[cs_ii][31:8]});
        
        // If the second half of the cs field is the inverse of the first then
        // sample the data
        wire rx_csf_err_free = rx_csf[63:32] == ~(rx_csf[31:0]);

        // If the data on this lane will be sampled, then indicate that the idle2
        // field was completely received to the CFG space.
        always @(posedge gt_pcs_clk) begin
          if (gt_pcs_rst_q) begin
            sample_csf_data       <= #TCQ 0;
            PPR_idle2_rcvd[cs_ii] <= #TCQ 0;
          end else begin
            if (sample_csf_data) begin
              sample_csf_data       <= #TCQ 0;
              PPR_idle2_rcvd[cs_ii] <= #TCQ 0;
            end else if (PPR_idle2_selected && cs_ctr_en_qqq && !cs_ctr_en_qq) begin
              sample_csf_data       <= #TCQ rx_csf_err_free;
              PPR_idle2_rcvd[cs_ii] <= #TCQ rx_csf_err_free;
            end
          end
        end 

        //*COVERAGE*
        // (cp_cs_start) : Cover all the valid combinations of the cs_start_q field
        // set illegal bins for bad values
        
        wire cs_aligned = cs_start[3] || cs_start_q[3]; // 4'b1000

        // Save the entire decoded CS field as it arrives to check of validity
        // of sampling its data.
        always @(posedge gt_pcs_clk) begin
          if (gt_pcs_rst_q) begin
            rx_csf <= #TCQ 0;
          end else begin
            // Select the data and decode it after the CS Field Marker completes
            // Aligned case contains all 8 bit on the same cycle
            // cs_ctr_en* should not be asserted if the field is interrupted or contains bit errors
            if (cs_ctr_en_q && cs_aligned) begin
              // Subtract 1 from the ctr to account for the second half of the csfm
              // Start filling on the LHS
              rx_csf[(8-(cs_ctr-1)-1)*8+:8] <= #TCQ decode_1000;

            // Mis-Aligned cases take an extra cycles to get all 4 cs field bytes
            end else if (cs_ctr_en_qq && !cs_aligned) begin
              // Subtract 2, one for the second half of the csfm and another for 
              // the extra cycle it takes to get the first full 32-bits of cs data
              case (cs_start_q)
                4'b0100: rx_csf[(8-(cs_ctr-2)-1)*8+:8] <= #TCQ decode_0100;
                4'b0010: rx_csf[(8-(cs_ctr-2)-1)*8+:8] <= #TCQ decode_0010;
                4'b0001: rx_csf[(8-(cs_ctr-2)-1)*8+:8] <= #TCQ decode_0001;
                default: rx_csf[(8-(cs_ctr-2)-1)*8+:8] <= #TCQ 8'bX;
              endcase

            //Clear this field whenever it is not being sampled.
            end else if (!rx_csf_err_free) begin
              rx_csf <= #TCQ 0;
            end
          end
        end

        // Sample the port width and lane number from the cs field only
        // if the CSFM doesnt contain an error.
        always @(posedge gt_pcs_clk) begin
          if (gt_pcs_rst_q) begin
            rx_port_width  <= #TCQ 0;
            rx_lane_number <= #TCQ 0;
          end else begin
            // Aligned case data is all available on the first cycle
            if (cs_ctr_en && !cs_ctr_en_q && cs_aligned &&
               (rx_data_exp[cs_ii][23:16] == ~rx_data_exp[cs_ii][7:0])) begin
              rx_port_width  <= #TCQ rx_data_exp[cs_ii][23:21];
              rx_lane_number <= #TCQ rx_data_exp[cs_ii][19:16];
            end 
            // Mis-aligned case
            else if (cs_ctr_en_q && !cs_ctr_en_qq && !cs_aligned) begin
               case (cs_start_q)
                4'b0100: begin
                  if (rx_data_exp_q[cs_ii][15:8] == ~rx_data_exp[cs_ii][31:24]) begin
                    rx_port_width  <= #TCQ rx_data_exp_q[cs_ii][15:13];
                    rx_lane_number <= #TCQ rx_data_exp_q[cs_ii][11:8];
                  end
                end
                4'b0010: begin
                  if (rx_data_exp_q[cs_ii][7:0] == ~rx_data_exp[cs_ii][23:16]) begin
                    rx_port_width  <= #TCQ rx_data_exp_q[cs_ii][7:5];
                    rx_lane_number <= #TCQ rx_data_exp_q[cs_ii][3:0];
                  end
                end
                4'b0001: begin
                  if (rx_data_exp[cs_ii][31:24] == ~rx_data_exp[cs_ii][15:8]) begin
                    rx_port_width  <= #TCQ rx_data_exp[cs_ii][31:29];
                    rx_lane_number <= #TCQ rx_data_exp[cs_ii][27:24];
                  end
                end
                default: begin
                  rx_port_width  <= #TCQ 3'bX;
                  rx_lane_number <= #TCQ 4'bX;
                end
              endcase
            end
          end
        end

        // Strip off the upper half on the rx_csf so we just have the non-inverted
        // data this way, when stripping off bits the bit index is intuitive 
        wire [31:0] rx_csf_validbits = rx_csf[63:32];

        // If the core is trained, dont sample the CS field for invalid
        // operating lanes even if there is one present
        wire valid_lane = !PPI_mode_1x || 
                          (PPI_mode_1x &&  PPI_rx_lane_r && (cs_ii == R)) ||
                          (PPI_mode_1x && !PPI_rx_lane_r && (cs_ii == 0));

        always @(posedge gt_pcs_clk) begin
          if (gt_pcs_rst_q) begin
            PPR_rx_port_width[cs_ii*3+:3]       <= #TCQ 0;
            PPR_rx_lane_number[cs_ii*4+:4]      <= #TCQ 0;
            PPR_receiver_trained[cs_ii]         <= #TCQ 0;
            PPR_gtrx_tap_p1_status[cs_ii*2+:2]  <= #TCQ 0;
            PPR_gtrx_tap_m1_status[cs_ii*2+:2]  <= #TCQ 0;
            PPR_rx_scram_en[cs_ii]              <= #TCQ 0;
            PPR_gtrx_cmd[cs_ii]                 <= #TCQ 0;
            PPR_gtrx_tap_m1_cmd[cs_ii*2+:2]     <= #TCQ 0;
            PPR_gtrx_tap_p1_cmd[cs_ii*2+:2]     <= #TCQ 0;
            PPR_gtrx_reset_emphasis[cs_ii]      <= #TCQ 0;
            PPR_gtrx_preset_emphasis[cs_ii]     <= #TCQ 0;
            PPR_gtrx_ack[cs_ii]                 <= #TCQ 0;
            PPR_gtrx_nack[cs_ii]                <= #TCQ 0;

          end else begin
            if (sample_csf_data && valid_lane) begin
              PPR_rx_port_width[cs_ii*3+:3]       <= #TCQ rx_port_width;
              PPR_rx_lane_number[cs_ii*4+:4]      <= #TCQ rx_lane_number;
              PPR_gtrx_cmd[cs_ii]                 <= #TCQ rx_csf_validbits[31];
              PPR_receiver_trained[cs_ii]         <= #TCQ rx_csf_validbits[29];
              PPR_rx_scram_en[cs_ii]              <= #TCQ rx_csf_validbits[28];              
              PPR_gtrx_tap_m1_status[cs_ii*2+:2]  <= #TCQ rx_csf_validbits[27:26];
              PPR_gtrx_tap_p1_status[cs_ii*2+:2]  <= #TCQ rx_csf_validbits[25:24];
              PPR_gtrx_tap_m1_cmd[cs_ii*2+:2]     <= #TCQ rx_csf_validbits[7:6];
              PPR_gtrx_tap_p1_cmd[cs_ii*2+:2]     <= #TCQ rx_csf_validbits[5:4];
              PPR_gtrx_reset_emphasis[cs_ii]      <= #TCQ rx_csf_validbits[3];
              PPR_gtrx_preset_emphasis[cs_ii]     <= #TCQ rx_csf_validbits[2];
              PPR_gtrx_ack[cs_ii]                 <= #TCQ rx_csf_validbits[1];
              PPR_gtrx_nack[cs_ii]                <= #TCQ rx_csf_validbits[0];
            end
          end
        end
      end //end for (cs_ii < LINK_WIDTH)

    end else begin : no_cs_decoder_gen
      //Tie off output signals to the PCFG if not in IDLE2 mode
      always @(posedge gt_pcs_clk) begin
        PPR_idle2_rcvd            <= #TCQ 0;
        PPR_receiver_trained      <= #TCQ 0;
        PPR_gtrx_tap_p1_status    <= #TCQ 0;
        PPR_gtrx_tap_m1_status    <= #TCQ 0;
        PPR_rx_scram_en           <= #TCQ 0;
        PPR_rx_port_width         <= #TCQ 0;
        PPR_rx_lane_number        <= #TCQ 0;
        PPR_gtrx_cmd              <= #TCQ 0;
        PPR_gtrx_tap_m1_cmd       <= #TCQ 0;
        PPR_gtrx_tap_p1_cmd       <= #TCQ 0;
        PPR_gtrx_reset_emphasis   <= #TCQ 0;
        PPR_gtrx_preset_emphasis  <= #TCQ 0;
        PPR_gtrx_ack              <= #TCQ 0;
        PPR_gtrx_nack             <= #TCQ 0;
      end
    end //if (!IDLE2)
  endgenerate
  // }}} Command and Status Decoder --------

  // {{{ + Descramblers + ------------------
  //Generate a descrambler for each lane
  //These are created outside the scope of the generate in order to assist
  //in coverage in the bind files.  This enables automatic binding and
  //eliminates the need for heirarchical references.
  reg   [GT_BYTES-1:0]    sync_check_reset  [LINK_WIDTH-1:0];
  wire  [16:0]            lfsr1_curr        [LINK_WIDTH-1:0];
  wire  [16:0]            lfsr2_curr        [LINK_WIDTH-1:0];
  wire  [16:0]            lfsr1_8           [LINK_WIDTH-1:0];
  reg   [GT_BYTES-1:0]    charisk_q         [LINK_WIDTH-1:0];
  reg   [GT_BYTES-1:0]    charisr_q         [LINK_WIDTH-1:0];
  reg   [GT_BYTES-1:0]    charism_q         [LINK_WIDTH-1:0];

  //For IDLE2 mode generate the logic to detect the CS Field of the idle2
  //sequence.
  genvar csb_ii;
  generate if (IDLE2) begin: cs_field_gen
    // {{{ CS Field Identification -----
    reg [1:0] master_lane;

    //CS Field counter
    //The cs field starts after two M's are detected. Use lane 0 as the 
    //master lane since they are all identical in the idle sequence
    //The charism wire is assigned in the scrambler generation blocks.
    //so we dont need duplicate logic here to assign it.
    
    //Figure out which lane to monitor as the master
    //If we are in 1x mode, use the lane with sync on it, otherwise just use
    //lane 0.
    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        master_lane <= #TCQ 0;
      end else begin
        master_lane <= #TCQ (PPI_mode_1x || (LINK_WIDTH == 1)) ? 
                              (PPI_lane_sync[0] ? 2'b0 : R) : 2'b0;
      end
    end

    //*ASSERTION*
    //(ap_cs_start): the start of the cs field is a one hot zero signal

    //*COVERPOINT*
    //(cp_csmarker_alignment): the CS field markers arrive in all alignment combinations

    //*COVERAGE*
    //(cp_cs_start_multiple_locations): See the cs field start with more than 4 M's, this is an 
    // error condition.

    assign cs_start_d[3] = &charism_q[master_lane];
    assign cs_start_d[2] = &charism_q[master_lane][2:0] &&  rx_charism_exp[master_lane][3];
    assign cs_start_d[1] = &charism_q[master_lane][1:0] && &rx_charism_exp[master_lane][3:2];
    assign cs_start_d[0] =  charism_q[master_lane][0]   && &rx_charism_exp[master_lane][3:1];

    // Protect against more than 4 /M/ characters starting the cs field. assume the last /M/ 
    // as the starting location
    always @* begin
      casex (cs_start_d)
        4'b0000: cs_start = 4'b0000;
        4'b1000: cs_start = 4'b1000;
        4'bx100: cs_start = 4'b0100;
        4'bxx10: cs_start = 4'b0010;
        4'bxxx1: cs_start = 4'b0001;
        default: cs_start = 4'bX;
      endcase
    end

    // Save the starting cs location to know what the current bytes alignment of the cs field is
    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        cs_start_q <= #TCQ 0;
      end else begin
        // As soon as enable asserts latch the start location
        if (cs_ctr_en && !cs_ctr_en_q) begin
          cs_start_q <= #TCQ cs_start;
        end
      end
    end

    // The cs field is interrupt whenever there is a K char seen. (this can
    // not be an M in which case its the csfield marker) 
    // If a bytes is interrupted, everything after it is too since that is no long 
    // the cs_field (this is needed to scrambler properly on an interrupt)
    assign cs_interrupt[3] = rx_chariskchar_exp[master_lane][3] && !rx_charism_exp[master_lane][3];
    assign cs_interrupt[2] = (rx_chariskchar_exp[master_lane][2] && !rx_charism_exp[master_lane][2]) || 
                             cs_interrupt[3];
    assign cs_interrupt[1] = (rx_chariskchar_exp[master_lane][1] && !rx_charism_exp[master_lane][1]) || 
                             cs_interrupt[2];
    assign cs_interrupt[0] = (rx_chariskchar_exp[master_lane][0] && !rx_charism_exp[master_lane][0]) || 
                             cs_interrupt[1];

    //*COVERAGE*
    //(cp_cs_interrupt): An cs field interrupt occurs in all valid combinations

    //*COVERAGE*
    //(cp_cs_interrupt_after_m): The cs field is interrupted after the 4 M's are detected

    //*COVERAGE*
    //(cp_cs_interrupt_after_marker): The cs field is interrupted after the entire cs field marker

    //*COVERAGE*
    //(cp_cs_interrupt_mid): The cs field is interrupted mid stream

    always @(*) begin
      // At the end of the cs_field, or if the csfield gets interrupted,
      // disable the counter
      if ((cs_ctr == CS_CYCLES-1) || |cs_interrupt) begin
        cs_ctr_en = 1'b0;
      end else if (|cs_start) begin
        cs_ctr_en = 1'b1;
      end else begin
        cs_ctr_en = cs_ctr_en_q;
      end
    end
        
    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        cs_ctr_en_q <= #TCQ 0;
      end else begin
        // Reset this at ctr-2 since this is what is used to figure out cs_field
        if ((cs_ctr == CS_CYCLES-2) || |cs_interrupt) begin
          cs_ctr_en_q <= #TCQ 0;
        end else begin
          cs_ctr_en_q <= #TCQ cs_ctr_en;
        end
      end
    end

    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        cs_ctr_en_qq <= #TCQ 0;
        cs_ctr_en_qqq <= #TCQ 0;
      end else begin
        cs_ctr_en_qq <= #TCQ cs_ctr_en_q;
        cs_ctr_en_qqq <= #TCQ cs_ctr_en_qq;
      end
    end

    //*ASSERTION*
    //(ap_cs_ctr_overcount): the cs_ctr does not count past CS_CYCLES
    
    //Count the number of cs field bytes
    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        cs_ctr <= #TCQ 0;
      end else begin
        if (cs_ctr_en) begin
          cs_ctr <= #TCQ cs_ctr + 1'b1;
        end else begin
          cs_ctr <= #TCQ 0;
        end
      end
    end

    //This is part of the cs field if the enable is asserted.  If it is
    //the first cycle, the bit in which the cs field started only asserts
    //If it is the last cycle, we know which bit is part of the cs field
    //by the number of bytes counted so far.
    for (csb_ii=0; csb_ii < GT_BYTES; csb_ii=csb_ii+1) begin: cs_field_gen
      assign cs_field[csb_ii] = (cs_ctr_en_q || cs_start[GT_BYTES-1:csb_ii]) && 
                                !cs_interrupt[csb_ii];
    end      
    //*COVERPOINT*
    //(cp_cs_field): the cs_field signal shows an offset cs field
    // }}} CS Field Identification -----
  end else begin: no_cs_field_gen
    assign cs_interrupt = 0;
    always @(posedge gt_pcs_clk) begin
      cs_ctr <= #TCQ 0;
    end
  end endgenerate

  //For IDLE2 cores, generate the logic to detect the command and status
  genvar dl_ii;   // descrambler lanes
  genvar dxor_ii; // descrambler xor
  genvar ll_ii;   // lfsr load
  genvar df_ii;   // descrambler fail
  genvar db_ii;   // descrambler bypass
  genvar dsl_ii;  // destripe lanes
  genvar dsb_ii;  // destripe bytes

  wire  [LINK_WIDTH-1:0]  load_by_lower_m;
  reg   [LINK_WIDTH-1:0]  load_by_upper_m;
  wire  [GT_BYTES-1:0]    sync_check_start    [LINK_WIDTH-1:0];
  reg   [GT_BYTES-1:0]    sync_check_stage1   [LINK_WIDTH-1:0];
  reg   [GT_BYTES-1:0]    sync_check_stage2   [LINK_WIDTH-1:0];

  generate if (IDLE2) begin: descrambler_gen
    //Generate a descrambler for each lane
    for (dl_ii=0; dl_ii < LINK_WIDTH; dl_ii=dl_ii+1) begin: descram_lane_gen
      //Declare Wires local to each scrambler
      wire                   load;
      wire                   shift16_on_load;
      wire  [GT_BYTES*8-1:0] descrambled_data;
      wire  [16:0]           load_data;
      wire  [16:0]           lfsr_load;
      reg   [GT_BYTES-1:0]   descram_fail;
      wire  [GT_BYTES-1:0]   bypass_descram;
      reg                    sync_failure;

      //*COVERPOINT*
      //(cp_charisr): Cover all interesting cases of charis R occur for IDLE2 only

      //*COVERPOINT*
      //(cp_charisk): Cover all interesting cases of charis R occur for IDLE2 only

      //*COVERPOINT*
      //(cp_charism): Cover all interesting cases of charis R occur for IDLE2 only

      //*COVERPOINT*
      //(cp_chariskchar): Cover all interesting combinations of charisk for IDLE2 only

      //Register char is R/K/M to be used in the descrambler sync checker
      //charism is accessed differenet since it is used elsewhere in this
      //file and declared outside the scope of the generate for loop.
      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          charisr_q[dl_ii] <= #TCQ 0;
          charisk_q[dl_ii] <= #TCQ 0;
          charism_q[dl_ii] <= #TCQ 0;
        end else begin
          charisr_q[dl_ii] <= #TCQ rx_charisr_exp[dl_ii];
          charisk_q[dl_ii] <= #TCQ rx_charisk_exp[dl_ii];
          charism_q[dl_ii] <= #TCQ rx_charism_exp[dl_ii];
        end
      end

      //Register the rx_data to know when to load the LFSR and
      //values to sample of the cs field
      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          rx_data_exp_q[dl_ii]         <= #TCQ 0;
          rx_chariskchar_exp_q[dl_ii]  <= #TCQ 0;
        end else begin
          rx_data_exp_q[dl_ii]         <= #TCQ rx_data_exp[dl_ii];
          rx_chariskchar_exp_q[dl_ii]  <= #TCQ rx_chariskchar_exp[dl_ii];
        end
      end

      // {{{ LFSR ------------------------

      // A load into the LFSR must occur whenever only one M character is seen. 
      // It should not load if the M is from the CS field
      // The load_by_.._m signals should assert on the cycle all 17 data bits to load are available.
      // M D D D | D 
      // X M D D | D D
      // X X M D | D D D
      // X X X M | D D D
      // Load by lower cant assert until it checks that the current data cycle is not part of the CS field
      // which occurs the cycle after an /M/ so this is not register
      // Load by upper knows wether it is in the cs field on the same cycle so it can be registered
      assign load_by_lower_m[dl_ii] = (!charism_q[dl_ii][2] && charism_q[dl_ii][1] && 
                                       !charism_q[dl_ii][0]) ||
                                      (!charism_q[dl_ii][1] && charism_q[dl_ii][0] && 
                                       !rx_charism_exp[dl_ii][3]);

      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          load_by_upper_m[dl_ii] <= #TCQ 0;
        end else begin
          load_by_upper_m[dl_ii] <= #TCQ (!charism_q[dl_ii][0] && rx_charism_exp[dl_ii][3] && 
                                          !rx_charism_exp[dl_ii][2]) ||
                                         (!rx_charism_exp[dl_ii][3] && rx_charism_exp[dl_ii][2] && 
                                          !rx_charism_exp[dl_ii][1]);
        end
      end

      //*COVERAGE*
      //(cp_load_by_upper_m): A scrambler load occurs from seeing an M on the upper two bytes

      //*COVERAGE*
      //(cp_load_by_lower_m): A scrambler load occurs from seeing an M on the lower two bytes

      // Based on the location of the /M/ grab 17 bits to load with
      assign load_data = load_by_upper_m[dl_ii] ? {rx_data_exp_q[dl_ii][15:0],rx_data_exp[dl_ii][31]} :
                                                  rx_data_exp[dl_ii][31:15];

      // A load occurs whenever an M is detected and this lane is out of sync
      assign load = (load_by_lower_m[dl_ii] || load_by_upper_m[dl_ii]) && ln_out_of_sync[dl_ii];

      // If the /M/ was detected on the upper bits we need to shift by 16 before loading
      // this is required since we need to use bytes from the previous cycle to load with
      // and it was shifted.
      assign shift16_on_load = load_by_upper_m[dl_ii] ?  1'b1 : 1'b0;

      // Reserve the incoming data since to load the LFSR with
      for (ll_ii=0; ll_ii < 17; ll_ii=ll_ii+1) begin: load_value_gen
        assign lfsr_load[16-ll_ii] = load_data[ll_ii];
      end //end for (ll_ii < 32)

      wire [2:0] r_count = rx_charisr_exp[dl_ii][0] + rx_charisr_exp[dl_ii][1] + 
                           rx_charisr_exp[dl_ii][2] + rx_charisr_exp[dl_ii][3];

      srio_gen2_v4_1_16_oplm_lfsr #(
        .TCQ          (TCQ),
        .LANE         (dl_ii),    
        .DESCRAMBLER  (1)
      ) oplm_lfsr1_rx_inst (   
        .gt_pcs_clk        (gt_pcs_clk),     
        .gt_pcs_rst_q      (gt_pcs_rst_q),
        .load              (load),
        .shift16_on_load   (shift16_on_load),
        .load_value        (lfsr_load),
        .r_count           (r_count),  
        .lfsr_curr         (lfsr1_curr[dl_ii]),
        .lfsr_8            (lfsr1_8[dl_ii]) 
      );
      srio_gen2_v4_1_16_oplm_lfsr #(
        .TCQ          (TCQ),
        .LANE         (dl_ii),    
        .DESCRAMBLER  (2)
      ) oplm_lfsr2_rx_inst (   
        .gt_pcs_clk        (gt_pcs_clk),
        .gt_pcs_rst_q      (gt_pcs_rst_q),
        .load              (load),
        .shift16_on_load   (shift16_on_load),
        .load_value        (lfsr_load),
        .r_count           (r_count),  
        .lfsr_curr         (lfsr2_curr[dl_ii]),
        .lfsr_8            () 
      );

      // }}} LFSR ------------------------

      // {{{ Descrambler Synchronization Checker
      // Look at the data stream for a K/M/R followed by data. When this occurs a sync check
      // should be performed on 4 bytes of data which is must results in D0.0's
      // This should not occur from any /M/ characters which starts the cs field
      assign sync_check_start[dl_ii][3] = (rx_charisk_exp[dl_ii][3] || rx_charism_exp[dl_ii][3] ||
                                           rx_charisr_exp[dl_ii][3]) && 
                                           !(|rx_chariskchar_exp[dl_ii][2:0]) && !charism_q[dl_ii][0]  && !(|cs_field);

      assign sync_check_start[dl_ii][2] = (rx_charisk_exp[dl_ii][2] || rx_charism_exp[dl_ii][2] ||
                                           rx_charisr_exp[dl_ii][2]) && 
                                           !(|rx_chariskchar_exp[dl_ii][1:0]) && !rx_charism_exp[dl_ii][3]  && !(|cs_field);
      assign sync_check_start[dl_ii][1] = (rx_charisk_exp[dl_ii][1] || rx_charism_exp[dl_ii][1] ||
                                           rx_charisr_exp[dl_ii][1]) && 
                                           !rx_chariskchar_exp[dl_ii][0] && !rx_charism_exp[dl_ii][2] && !(|cs_field);

      assign sync_check_start[dl_ii][0] = (rx_charisk_exp[dl_ii][0] || rx_charism_exp[dl_ii][0] ||
                                           rx_charisr_exp[dl_ii][0]) && !rx_charism_exp[dl_ii][1]  && !(|cs_field);


      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          sync_check_reset[dl_ii]   <= #TCQ 0; 
          sync_check_stage1[dl_ii]  <= #TCQ 0;
          sync_check_stage2[dl_ii]  <= #TCQ 0;
        end else begin
          // If we are already out of sync, or reloading dont perform new sync
          // checks
          if (|ln_out_of_sync || load) begin
            sync_check_reset[dl_ii]   <= #TCQ 0;
            sync_check_stage1[dl_ii]  <= #TCQ 0;
            sync_check_stage2[dl_ii]  <= #TCQ 0;

          end else begin
            sync_check_reset[dl_ii]   <= #TCQ rx_chariskchar_exp[dl_ii] | rx_invalid_exp[dl_ii];
            sync_check_stage1[dl_ii]  <= #TCQ sync_check_start[dl_ii];
            sync_check_stage2[dl_ii]  <= #TCQ sync_check_stage1[dl_ii];
          end
        end
      end

      //*ASSERTION*
      // (ap_sync_check_in_cs): A sync check is not issued while in the cs field
      
      //*COVERPOINT*
      //(cp_sync_check_interrupt_start): A K character interrupts a sync check start
      //(cp_sync_check_interrupt_stage1): A K character interrupts a sync check in stage1
      //(cp_sync_check_interrupt_stage2): A K character interrupts a sync check in stage2
      
      // Register this data for the check data
      for (df_ii=0; df_ii < GT_BYTES; df_ii=df_ii+1) begin: descram_fail_gen
        always @(posedge gt_pcs_clk) begin
          if (gt_pcs_rst_q) begin
            descram_fail[df_ii] <= #TCQ 0;
          end else begin
            descram_fail[df_ii] <= #TCQ !rx_chariskchar_exp[dl_ii][df_ii] && 
                                        |descrambled_data[df_ii*8+:8];
          end
        end
      end //end for (df_ii < GT_BYTES)

      //A sync check has failed if there is not a K character and the data
      //did not come out to be 0's
      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          sync_failure  <= #TCQ 0;

        end else begin
          // If we are loading a new descrambler value dont fail further
          // checks until the next sync check starts
          if (load) begin
            sync_failure  <= #TCQ 0;

          end else if (|sync_check_stage1[dl_ii]) begin
            casex (sync_check_stage1[dl_ii]) 
              4'b1xxx: sync_failure <= #TCQ |descram_fail[2:0] && !(|sync_check_reset[dl_ii][1:0]);
              4'b01xx: sync_failure <= #TCQ |descram_fail[1:0] && !(|sync_check_reset[dl_ii][1:0]);
              4'b001x: sync_failure <= #TCQ  descram_fail[0]   && !sync_check_reset[dl_ii][0];
              4'b0001: sync_failure <= #TCQ 0; //check all 4 bytes in stage2 on next cycle
              default: sync_failure <= #TCQ 1'bX;
            endcase

          end else if (sync_check_stage2[dl_ii]) begin
            casex (sync_check_stage2[dl_ii]) 
              4'b1xxx: sync_failure <= #TCQ descram_fail[3]    && !sync_check_reset[dl_ii][3];
              4'b01xx: sync_failure <= #TCQ |descram_fail[3:2] && !(|sync_check_reset[dl_ii][3:2]);
              4'b001x: sync_failure <= #TCQ |descram_fail[3:1] && !(|sync_check_reset[dl_ii][3:1]);
              4'b0001: sync_failure <= #TCQ |descram_fail      && !(|sync_check_reset[dl_ii]);
              default: sync_failure <= #TCQ 1'bX;
            endcase
          end else begin
            sync_failure <= #TCQ 0;
          end
        end 
      end //end always

      //Drive the descrambler out of sync signal for this descrambler.  If 
      //any sync check does not pass, the descrambler is out of sync.
      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          ln_out_of_sync[dl_ii] <= #TCQ 1;
        end else begin
          if (load || (SCRAM == 0)) begin
            ln_out_of_sync[dl_ii] <= #TCQ 0;

          end else if (sync_failure) begin
            ln_out_of_sync[dl_ii] <= #TCQ 1;
          end
        end
      end

      //*COVERAGE*
      // (cp_ln_out_of_sync): Cover all combination of lanes of out sync

      // }}} Descrambler Synchronization Checker

      //When scrambing the data the lfsr_scram uses a 1:17 methodology to
      //match the spec for bit "16" needs to be XORed with bit "15" of the
      //data since bit 15 will go out first.
      //Shifting matches these cases (these are boiled down from looking at K/R/M locations with 1-5 Rs):
      //  A:  RMxx  (sh8)
      //  B:  RRMx  (sh16)
      //  C:  KRMx  (sh8)
      wire [31:0] lfsr_curr = (r_count == 1 && (rx_charisr_exp[dl_ii][3] || rx_charisr_exp[dl_ii][2]))  ?
                               {lfsr1_8[dl_ii][15:0], lfsr1_curr[dl_ii][15:0]} :
                              (r_count == 2 && rx_charisr_exp[dl_ii][2])  ?
                               {lfsr1_curr[dl_ii][15:0], lfsr1_curr[dl_ii][15:0]} :
                               {lfsr2_curr[dl_ii][15:0], lfsr1_curr[dl_ii][15:0]};

      for (dxor_ii=0; dxor_ii < 32; dxor_ii=dxor_ii+1) begin: descrambled_data_xor_gen
        assign descrambled_data[31-dxor_ii] = rx_data_exp[dl_ii][31-dxor_ii] ^ lfsr_curr[dxor_ii];
      end

      //Check data bytes for descrambling. Descramble if:
      //1. Scrambling is not allowed in the system
      //2. it is not a K character
      //3. is is not the cs field
      //4. it is not the idle field and PC_scram_disable is set
      for (db_ii=0; db_ii < GT_BYTES; db_ii=db_ii+1) begin : descram_gen
        assign bypass_descram[db_ii] = !PPR_idle2_selected || (SCRAM == 0) || cs_field[db_ii] ||
                                       rx_chariskchar_exp[dl_ii][db_ii] ||
                                       (PC_scram_disable && (descrambled_data[db_ii*8+:8] != 0));

        always @(posedge gt_pcs_clk) begin
          if (gt_pcs_rst_q) begin
            descram[dl_ii][db_ii*8+:8] <= #TCQ 0;
          end else begin
            descram[dl_ii][db_ii*8+:8] <= #TCQ bypass_descram[db_ii] ? rx_data_exp[dl_ii][db_ii*8+:8] :
                                                                       descrambled_data[db_ii*8+:8];
          end
        end
      end //end for (db_ii < GT_BYTES)

      //Pass on K characters and any GT errors
      always @(posedge gt_pcs_clk) begin
        if (gt_pcs_rst_q) begin
          descram_isk[dl_ii]     <= #TCQ 0;
          descram_invalid[dl_ii] <= #TCQ 0;
          descram_pd_sc[dl_ii]   <= #TCQ 0;
        end else begin
          descram_isk[dl_ii]     <= #TCQ rx_chariskchar_exp[dl_ii];
          descram_invalid[dl_ii] <= #TCQ rx_invalid_exp[dl_ii];
          descram_pd_sc[dl_ii]   <= #TCQ rx_charispdsc_exp[dl_ii];
        end
      end
    end //end for (dl_ii < LANE_WIDTH)

    //Create of out of sync signal to pass to the OLLM. If any descrambler
    //is out of sync then drive this signal high. Only indicate out of sync when
    //operating in idle2 mode.
    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        gt_out_of_sync <= #TCQ 1;
      end else begin
        if (!PPR_idle2_selected) begin
          gt_out_of_sync <= #TCQ 0;

        end else begin
          if (PPI_mode_1x) begin
            gt_out_of_sync <= #TCQ (PPI_rx_lane_r) ? ln_out_of_sync[R] : ln_out_of_sync[0];
          end else begin
            gt_out_of_sync <= #TCQ |ln_out_of_sync;
          end
        end
      end
    end

    //*ASSERTION*
    //(ap_outofsync): If any lane is out of sync then the out of sync signal must assert
    //(ap_outofsync): on the next cycle.

  end else begin: no_descramer_gen
    always @(posedge gt_pcs_clk) begin
      gt_out_of_sync  <= #TCQ 0;
      load_by_upper_m <= #TCQ 0;
    end

    //Tie off these signals for the bind files
    wire   start_cs         = 0;
    assign load_by_lower_m  = 0;

    //Generate a tied off signals per lane
    for (dl_ii=0; dl_ii < LINK_WIDTH; dl_ii=dl_ii+1) begin: nodescram_lane_gen
      assign sync_check_start[dl_ii] = 0;
      always @(posedge gt_pcs_clk) begin
        sync_check_reset[dl_ii]  <= #TCQ 0;
        sync_check_stage1[dl_ii]  <= #TCQ 0;
        sync_check_stage2[dl_ii]  <= #TCQ 0;
      end
    end
  end endgenerate //end if (IDLE2) for descrambler generation
  // }}} + Descramblers + ------------------

  // {{{ Destriping ------------------------
  generate
  for (dsb_ii=0; dsb_ii < GT_BYTES; dsb_ii=dsb_ii+1) begin: destripe_bytes_gen
    for (dsl_ii=0; dsl_ii < LINK_WIDTH; dsl_ii=dsl_ii+1) begin: destripe_gen_gen
      assign destripe_gen[((LINK_WIDTH*8*dsb_ii)+(dsl_ii*8))+:8] = (PPR_idle2_selected) ? 
                                                                   descram[LINK_WIDTH-1-dsl_ii][dsb_ii*8+:8] :
                                                                   rx_data_exp[LINK_WIDTH-1-dsl_ii][dsb_ii*8+:8];
      assign destripe_isk_gen[(LINK_WIDTH*dsb_ii+dsl_ii)]        = (PPR_idle2_selected) ? 
                                                                   descram_isk[LINK_WIDTH-1-dsl_ii][dsb_ii] :
                                                                   rx_chariskchar_exp[LINK_WIDTH-1-dsl_ii][dsb_ii];
      assign destripe_invalid_gen[(LINK_WIDTH*dsb_ii+dsl_ii)]    = (PPR_idle2_selected) ? 
                                                                   descram_invalid[LINK_WIDTH-1-dsl_ii][dsb_ii] :
                                                                   rx_invalid_exp[LINK_WIDTH-1-dsl_ii][dsb_ii];
      assign destripe_pdsc_gen[(LINK_WIDTH*dsb_ii+dsl_ii)]       = (PPR_idle2_selected) ? 
                                                                   descram_pd_sc[LINK_WIDTH-1-dsl_ii][dsb_ii] :
                                                                   rx_charispdsc_exp[LINK_WIDTH-1-dsl_ii][dsb_ii];
    end
  end
  endgenerate

  always @(posedge gt_pcs_clk) begin
    // No need to reset the data 
    if (gt_pcs_rst_q) begin
      destripe_invalid <= #TCQ 1;
      destripe_pdsc    <= #TCQ 0;

    //For 1x or trained cores, select either lane 0 or the redundancy lane R
    //based on the PPI_rx_lane_r signal from the initialization state machines.
    end else if (PPI_mode_1x) begin
      if (PPI_rx_lane_r) begin
        destripe          <= #TCQ (PPR_idle2_selected) ? descram[R]         : rx_data_exp[R];
        destripe_isk      <= #TCQ (PPR_idle2_selected) ? descram_isk[R]     : rx_chariskchar_exp[R];
        destripe_invalid  <= #TCQ (PPR_idle2_selected) ? descram_invalid[R] : rx_invalid_exp[R];
        destripe_pdsc     <= #TCQ (PPR_idle2_selected) ? descram_pd_sc[R]   : rx_charispdsc_exp[R];
      end else begin
        destripe          <= #TCQ (PPR_idle2_selected) ? descram[0]         : rx_data_exp[0];
        destripe_isk      <= #TCQ (PPR_idle2_selected) ? descram_isk[0]     : rx_chariskchar_exp[0];
        destripe_invalid  <= #TCQ (PPR_idle2_selected) ? descram_invalid[0] : rx_invalid_exp[0];
        destripe_pdsc     <= #TCQ (PPR_idle2_selected) ? descram_pd_sc[0]   : rx_charispdsc_exp[0];
      end
    end else begin 
      destripe          <= #TCQ destripe_gen;
      destripe_isk      <= #TCQ destripe_isk_gen;
      destripe_invalid  <= #TCQ destripe_invalid_gen;
      destripe_pdsc     <= #TCQ destripe_pdsc_gen;
    end  
  end

  //*COVERAGE*
  //(cp_destripe_pdsc): Cover all the interesting combinations of a PD/SC detection for 
  // long control symbols

  //*COVERAGE*
  //(cp_destripe_pdsc_short_cs): Cover all the interesting combinations of a PD/SC detection
  // for short control symbols
  // }}} Destriping ------------------------

  // {{{ Byte Alignment -------------------------
  // Register all incoming destriped signals in order to shift alignment as needed
  // and align pd/sc characters to word boundaries
  always @(posedge gt_pcs_clk) begin
    // No need to reset the data
    if (gt_pcs_rst_q) begin
      destripe_invalid_q  <= #TCQ 1;
    end else begin
      destripe_q          <= #TCQ destripe;
      destripe_isk_q      <= #TCQ destripe_isk;
      destripe_invalid_q  <= #TCQ destripe_invalid;
      destripe_pdsc_q     <= #TCQ destripe_pdsc[3:0];
    end
  end

  // Montior for the start of a control symbol so realignment
  // does not occur on the end of a long control symbol
  // It is the end of the control symbol one cycle later if we are in alignment
  // all other alignment scenarios take two cycles to complete a control symbol
  // after the start is seen
  wire csymbol_end_1x    = (|destripe_pdsc && destripe_pdsc[aligned_end_idx_1x]) ||
                           (!(|destripe_pdsc) && byte_alignment == 4'b1000 && csymbol_toggle_q) ||
                           (!(|destripe_pdsc) && byte_alignment != 4'b1000 && csymbol_toggle_qq);
  wire csymbol_start_1x  = |destripe_pdsc &&
                           (csymbol_monitor || destripe_pdsc[aligned_start_idx_1x]);

  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      csymbol_monitor <= #TCQ 1;
    end else begin
      if (!IDLE2 || !PPI_port_initialized) begin
        csymbol_monitor <= #TCQ 1;

      end else if (PPI_mode_1x) begin
        if (csymbol_start_1x && PPR_idle2_selected) begin
          csymbol_monitor <= #TCQ 0;
        end else if (csymbol_end_1x && !csymbol_start_1x && PPR_idle2_selected) begin
          csymbol_monitor <= #TCQ 1;
        end

      end else if (LINK_WIDTH == 2 && PPR_idle2_selected) begin
        if (csymbol_start_2x && !csymbol_end_2x) begin
          csymbol_monitor <= #TCQ 0;
        end else if (csymbol_end_2x && !csymbol_start_2x) begin
          csymbol_monitor <= #TCQ 1;
        end
      end
    end
  end

  // When a stream of non-k characters occurs reset the start detect signal
  // this is needed for bad delimiters on control symbols.
  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      csymbol_toggle_q   <= #TCQ 0;
      csymbol_toggle_qq  <= #TCQ 0;
    end else begin
      csymbol_toggle_q   <= #TCQ (PPI_mode_1x) ? csymbol_start_1x : csymbol_start_2x;
      csymbol_toggle_qq  <= #TCQ csymbol_toggle_q;
    end
  end

  // The PD/SC character on byte 3 otherwise it is out of alignment for a x1 core
  always @* begin
    case (byte_alignment_q)
      4'b1000: aligned_start_idx_1x = 3;
      4'b0100: aligned_start_idx_1x = 2;
      4'b0010: aligned_start_idx_1x = 1;
      4'b0001: aligned_start_idx_1x = 0;
      default: aligned_start_idx_1x = 2'bX;
    endcase
  end

  always @* begin
    case (byte_alignment_q)
      4'b1000: aligned_end_idx_1x = 0;
      4'b0100: aligned_end_idx_1x = 3;
      4'b0010: aligned_end_idx_1x = 2;
      4'b0001: aligned_end_idx_1x = 1;
      default: aligned_end_idx_1x = 2'bX;
    endcase
  end

  assign correct_byte_alignment_1x = destripe_pdsc[aligned_start_idx_1x];

  // Based on the link width the alignment requirements change with the link width
  generate if (LINK_WIDTH == 1) begin: correct_byte_alignment_x1_gen
    assign correct_byte_alignment = correct_byte_alignment_1x;
    assign realign                = destripe_pdsc;
    assign valid_realign          = 1'b1;

  end else if (LINK_WIDTH == 2) begin: correct_byte_alignment_x2_gen
    reg aligned_end_idx_2x_q;

    always @* begin
      case (byte_alignment_q)
        4'b1000: aligned_start_idx_2x = 7;
        4'b0100: aligned_start_idx_2x = 6;
        4'b0010: aligned_start_idx_2x = 5;
        4'b0001: aligned_start_idx_2x = 4;
        default: aligned_start_idx_2x = 2'bX;
      endcase
    end

    always @(posedge gt_pcs_clk) begin
      if (csymbol_start_2x && !csymbol_end_2x) begin
        casex (destripe_pdsc)
          8'b1xxx_xxxx: aligned_end_idx_2x = 0;
          8'b01xx_xxxx: aligned_end_idx_2x = 7;
          8'b001x_xxxx: aligned_end_idx_2x = 6;
          8'b0001_xxxx: aligned_end_idx_2x = 5;
          8'b0000_1xxx: aligned_end_idx_2x = 4;
          8'b0000_01xx: aligned_end_idx_2x = 3;
          8'b0000_001x: aligned_end_idx_2x = 2;
          8'b0000_0001: aligned_end_idx_2x = 1;
          8'b0000_0000: aligned_end_idx_2x = aligned_end_idx_2x_q;
        default: aligned_end_idx_2x = 2'bX;
        endcase
      end
    end

    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        aligned_end_idx_2x_q <= #TCQ 0;
      end else begin
        aligned_end_idx_2x_q <= #TCQ aligned_end_idx_2x;
      end
    end

    assign csymbol_end_2x   = (|destripe_pdsc && !csymbol_monitor &&
                               (destripe_pdsc[aligned_end_idx_2x] || destripe_pdsc[aligned_end_idx_2x_lower])) ||
                              (byte_alignment == 4'b1000) && (destripe_pdsc[7]) ||
                              (!(|destripe_pdsc) && csymbol_toggle_q);
    assign csymbol_start_2x = |destripe_pdsc &&
                               (csymbol_monitor ||
                                destripe_pdsc[aligned_start_idx_2x_lower] ||
                                destripe_pdsc[aligned_start_idx_2x]);

    // If the starting index is 1000 or 0100 then there is an alternate alignment possible
    // otherwise there is not. This is because this is only checked on the starting delimiter.
    // This logic is only for long control symbols. For short, it is always re-aligning
    assign aligned_start_idx_2x_lower = (byte_alignment_q > 1) ? aligned_start_idx_2x-4 : aligned_start_idx_2x;
    assign aligned_end_idx_2x_lower   = (byte_alignment_q > 1) ? aligned_end_idx_2x-4 : aligned_end_idx_2x;

    assign correct_byte_alignment = (PPI_mode_1x) ? correct_byte_alignment_1x :
                                                    (destripe_pdsc[aligned_start_idx_2x_lower] ||
                                                     destripe_pdsc[aligned_start_idx_2x]) &&
                                                    (!multiple_alignments);

    assign realign = (PPI_mode_1x) ? destripe_pdsc[3:0] :
                                     (destripe_pdsc[7:4] | destripe_pdsc[3:0]);

    // In x1 any realign is allowed, in x2 mode dont realign if the pd/sc is on an invalid start lane
    assign valid_realign = (PPI_mode_1x) ? 1'b1 : destripe_pdsc[7] || destripe_pdsc[5] ||
                                                  destripe_pdsc[3] || destripe_pdsc[1];

  end else if (LINK_WIDTH == 4) begin: correct_byte_alignment_x4_genbegin
    // x4 cores are always in alignment unless its trained
    assign correct_byte_alignment = (PPI_mode_1x) ? correct_byte_alignment_1x : 1'b1;

    assign realign = (PPI_mode_1x) ? destripe_pdsc[3:0] : 4'b1000;

    // In x1 any realign is allowed, in x4 mode nothing should cause a realign
    assign valid_realign = (PPI_mode_1x) ? 1'b1 : 1'b0;
  end endgenerate

  //*COVERAGE*
  //(cp_byte_alignment): Cover all valid combinations of the byte alignment

  //*CROSS*
  //(cr_aligment_lw): cross all the byte_alignments with a x1 and x1 link width

  // If a delimiter is detected, check if the byte alignment is correct. If
  // the alignment check fail toggle the alignment to the other mode
  wire realign_allowed    = |realign && csymbol_monitor && valid_realign;
  wire new_byte_alignment = realign_allowed && !correct_byte_alignment;

  always @(*) begin
    if (new_byte_alignment) begin
      if (PPR_idle2_selected) begin
        casex (realign)
          4'b1xxx: byte_alignment = 4'b1000;
          4'b01xx: byte_alignment = 4'b0100;
          4'b001x: byte_alignment = 4'b0010;
          4'b0001: byte_alignment = 4'b0001;
          default: byte_alignment = 4'bx;
        endcase
      end else begin
        casex (realign)
          4'b1000: byte_alignment = 4'b1000;
          4'bx100: byte_alignment = 4'b0100;
          4'bxx10: byte_alignment = 4'b0010;
          4'bxxx1: byte_alignment = 4'b0001;
          default: byte_alignment = 4'bx;
        endcase
      end
    end else begin
      byte_alignment = byte_alignment_q;
    end
  end

  //latch the byte_alignment signal
  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      // Reset in an assumed aligned state
      byte_alignment_q  <= #TCQ 4'b1000;
      realign_allowed_q <= #TCQ 0;
      new_byte_alignment_q <= #TCQ 0;
    end else begin
      byte_alignment_q  <= #TCQ byte_alignment;
      realign_allowed_q <= #TCQ realign_allowed;
      new_byte_alignment_q <= #TCQ new_byte_alignment;
    end
  end

  // For a x1 core, data that realigns can have idles less than a cycle (ie
  // 3 bytes, while a cycle is 4 bytes) so shifting for alignment may result
  // in idle sequence errors. In this case, when we realign, insert idles
  // which will never result in an error to avoid rogue PNAs from the ollm rx
  wire [31:0] pad     = (PPR_idle2_selected) ? {D0_0,D0_0,D0_0,D0_0} : {R_CHAR,R_CHAR,R_CHAR,R_CHAR};
  wire [3:0]  pad_isk = (PPR_idle2_selected) ? 4'b0000 : 4'b1111;

  //*COVERAGE*
  //(cp_realign_x2):  See all the possible realignments on a x2
  //*ASSERTION*
  //(ap_realign_x4): A realign can not occur on a x4 link
  assign multiple_alignments = ((realign[3] + realign[2] + realign[1] + realign[0]) > 1) &&
                               !PPR_idle2_selected;

  always @* begin
    casex (realign)
      4'b1xxx: upper_byte_alignment = 4'b1000;
      4'b01xx: upper_byte_alignment = 4'b0100;
      4'b001x: upper_byte_alignment = 4'b0010;
      4'b0001: upper_byte_alignment = 4'b0001;
      default: upper_byte_alignment = 4'bx;
    endcase
  end

  //*ASSERTION*
  //(ap_multiple_alignments_x4): multiple_alignments can not assert on a x4 core


  // If the link is operating in x2 mode, we need to align differently since stripping does not allow us to use
  // the store/flush logic (only applies for each lane independently, but lane1 doesnt have pd/sc indicators to do this with).
  // This is occur when back2back control symbols are received and the alignment shifts left.
  wire rhs_b2b_cs = |destripe_pdsc_q[3:0] && |destripe_pdsc[3:0];
  wire left_shift = (destripe_pdsc_q[3:0] < destripe_pdsc[3:0]);
  wire shift_align_b2b_cs = rhs_b2b_cs && left_shift && new_byte_alignment;

  reg [31:0] realign_bytes;
  reg [3:0]  realign_isk;
  reg [3:0]  realign_invalid;

  always @* begin
    if (shift_align_b2b_cs) begin
      realign_bytes   = {destripe_q[0+:16], destripe[DATA_WIDTH-16+:16]};
      realign_isk     = {destripe_isk_q[0+:2], destripe_isk[CHARIS_WIDTH-2+:2]};
      realign_invalid = {destripe_invalid_q[0+:2], destripe_invalid[CHARIS_WIDTH-2+:2]};
    end else if (new_byte_alignment) begin
      realign_bytes   = pad[31:0];
      realign_isk     = pad_isk[3:0];
      realign_invalid = 4'b000;
    end else begin
      realign_bytes   = destripe_q[0+:31];
      realign_isk     = destripe_isk_q[0+:4];
      realign_invalid = destripe_invalid_q[0+:4];
    end
  end

  // Store bytes when the alignment mode switches
  wire flush_stored = new_byte_alignment && (byte_alignment > byte_alignment_q);

  //*COVERAGE*
  //(cr_flush_alignments): See a flush occur on all the possible alignments

  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      flush_stored_q <= #TCQ 0;
    end else begin
      flush_stored_q <= #TCQ flush_stored;
    end
  end

  wire [31:0] stored_bytes         = locked_bytes[1] ?
                                      {byte3_stored[7:0], byte2_stored[7:0], byte1_stored[7:0], destripe_q[7:0]} :
                                     locked_bytes[2] ?
                                      {byte3_stored[7:0], byte2_stored[7:0], destripe_q[15:0]} :
                                      {byte3_stored[7:0], destripe_q[23:0]};

  wire [3:0] stored_bytes_isk      = locked_bytes[1] ?
                                      {byte3_stored[8], byte2_stored[8], byte1_stored[8], destripe_isk_q[0]} :
                                     locked_bytes[2] ?
                                      {byte3_stored[8], byte2_stored[8], destripe_isk_q[1:0]} :
                                      {byte3_stored[8], destripe_isk_q[2:0]};

  wire [3:0] stored_bytes_invalid  = locked_bytes[1] ?
                                      {byte3_stored[9], byte2_stored[9], byte1_stored[9], destripe_invalid_q[0]} :
                                     locked_bytes[2] ?
                                      {byte3_stored[9], byte2_stored[9], destripe_invalid_q[1:0]} :
                                      {byte3_stored[9], destripe_invalid_q[2:0]};

  //*COVERAGE*
  // (cp_locked_bytes) : cover all the possible values of locked bytes

  //*COVERAGE*
  //(cr_locked_X_flush): See a flush on all the different locked cases

  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      locked_bytes <= #TCQ 0;
    end else if (new_byte_alignment) begin
      // Lock the necessary registers with their stored data until a flush
      // should occur
      case (byte_alignment)
        4'b1000: begin
          if (flush_stored) begin
            locked_bytes <= #TCQ 4'b0000;
          end else begin
            locked_bytes <= #TCQ ~locked_bytes[3];
          end
          locked_bytes <= #TCQ 0;
        end
        4'b0100: begin
          if (flush_stored) begin
            locked_bytes <= #TCQ 4'b1000;
          end else begin
            locked_bytes[3] <= #TCQ ~locked_bytes[3];
          end
          // Lock data from byte 3
          if (flush_stored || ~locked_bytes[3]) begin
            byte3_stored <= #TCQ {destripe_invalid[3],destripe_isk[3],destripe[31:24]};
          end
        end
        4'b0010: begin
          if (flush_stored) begin
            locked_bytes <= #TCQ 4'b1100;
          end else begin
            locked_bytes[3:2] <= #TCQ {2{~locked_bytes[2]}};
          end
          // Lock data from byte 3
          if (flush_stored || ~locked_bytes[3]) begin
            byte3_stored <= #TCQ {destripe_invalid[3],destripe_isk[3],destripe[31:24]};
          end
          // Lock data from byte 2
          if (flush_stored || ~locked_bytes[2]) begin
            byte2_stored <= #TCQ {destripe_invalid[2],destripe_isk[2],destripe[23:16]};
          end
        end
        4'b0001: begin
          if (flush_stored) begin
            locked_bytes <= #TCQ 4'b1110;
          end else begin
            locked_bytes[3:1] <= #TCQ {3{~locked_bytes[1]}};
          end
          // Lock data from byte 3
          if (flush_stored || ~locked_bytes[3]) begin
            byte3_stored <= #TCQ {destripe_invalid[3],destripe_isk[3],destripe[31:24]};
          end
          // Lock data from byte 2
          if (flush_stored || ~locked_bytes[2]) begin
            byte2_stored <= #TCQ {destripe_invalid[2],destripe_isk[2],destripe[23:16]};
          end
          // Lock data from byte 1
          if (flush_stored || ~locked_bytes[1]) begin
            byte1_stored <= #TCQ {destripe_invalid[1],destripe_isk[1],destripe[15:8]};
          end
        end
        default: locked_bytes <= #TCQ 4'bX;
      endcase
    end
  end

  // If the previous cycles was allowed to realign (meaning a PD/SC was seen), this cycle should use the
  // last value of the alignment otherwise that cycle will propigate out with a new alignment which is not
  // what we want.
  wire [3:0] byte_alignment_nx_d = (multiple_alignments) ? upper_byte_alignment : byte_alignment;

  //Set the rx data and sideband signals based on the alignment detected.
  //Invert the invalid signal to create a valid signal.  valid indicates that
  //there were not gt errors detected.
  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      // Only reset the control bits
      gt_rx_valid    <= #TCQ 0;
    end else begin
      if (PPI_mode_1x && !PPR_idle2_selected) begin
        case (byte_alignment_q)
        4'b1000: begin
          gt_rx_data     <= #TCQ (flush_stored) ? //stored_bytes      
                                   	                          // CR 824966, when the flush occurs there is no point in keeping old data and char bytes
	                                          32'hfdfdfdfd :  // /R/ bytes are chosen as clock compensation bytes
						  destripe_q;
          gt_rx_charisk  <= #TCQ (flush_stored) ? //stored_bytes_isk  
	                                          4'hf :          // CR 824966, all bytes are idle bytes, so all char bits are 1
						  destripe_isk_q;
          gt_rx_valid    <= #TCQ (flush_stored) ? ~stored_bytes_isk : ~destripe_invalid_q;
        end
        4'b0100: begin
          gt_rx_data    <= #TCQ (flush_stored) ? //stored_bytes :
                                                 32'hfdfdfdfd :   // CR 824966, when the flush occurs there is no point in keeping old data and char bytes
                                                 {destripe_q[0+:24], destripe[24+:32-24]};
          gt_rx_charisk <= #TCQ (flush_stored) ? //stored_bytes_isk :
	                                         4'hf :           // CR 824966, all bytes are idle bytes, so all char bits are 1
                                                 {destripe_isk_q[0+:3], destripe_isk[3+:4-3]};
          gt_rx_valid   <= #TCQ (flush_stored) ? ~stored_bytes_isk :
                                                 {~destripe_invalid_q[0+:3], ~destripe_invalid[3+:4-3]};
        end
        4'b0010: begin
          gt_rx_data    <= #TCQ (flush_stored) ? //stored_bytes :
	                                         32'hfdfdfdfd :   // CR 824966, when the flush occurs there is no point in keeping old data and char bytes
                                                 {destripe_q[0+:16], destripe[16+:32-16]};
          gt_rx_charisk <= #TCQ (flush_stored) ? //stored_bytes_isk :
	                                         4'hf :           // CR 824966, all bytes are idle bytes, so all char bits are 1
                                                 {destripe_isk_q[0+:2], destripe_isk[2+:4-2]};
          gt_rx_valid   <= #TCQ (flush_stored) ? ~stored_bytes_isk :
                                                 {~destripe_invalid_q[0+:2], ~destripe_invalid[2+:4-2]};
        end
        4'b0001: begin
          gt_rx_data    <= #TCQ (flush_stored) ? //stored_bytes :
	                                         32'hfdfdfdfd :   // CR 824966, when the flush occurs there is no point in keeping old data and char bytes
                                                 {destripe_q[0+:8], destripe[8+:32-8]};
          gt_rx_charisk <= #TCQ (flush_stored) ? //stored_bytes_isk :
	                                         4'hf :           // CR 824966, all bytes are idle bytes, so all char bits are 1
                                                 {destripe_isk_q[0+:1], destripe_isk[1+:4-1]};
          gt_rx_valid   <= #TCQ (flush_stored) ? ~stored_bytes_isk :
                                                 {~destripe_invalid_q[0+:1], ~destripe_invalid[1+:4-1]};
        end
        default: begin
          gt_rx_data    <= #TCQ {DATA_WIDTH{1'bX}};
          gt_rx_charisk <= #TCQ {CHARIS_WIDTH{1'bX}};
          gt_rx_valid   <= #TCQ {CHARIS_WIDTH{1'bX}};
        end
        endcase
        end else if (PPI_mode_1x && PPR_idle2_selected) begin
        case (byte_alignment_1x_d) 
        7'b0000001: begin // pass as is
                   gt_rx_data     <= #TCQ destripe;
                   gt_rx_charisk  <= #TCQ destripe_isk;
                   gt_rx_valid    <= #TCQ ~destripe_invalid;
                 end

        7'b0000010: begin // ONE_BIT_SHIFT
                  gt_rx_data     <= #TCQ {//destripe[63:32],
                                          destripe_q[7:0],
                                          destripe[31:8]
                                          };
                  gt_rx_charisk  <= #TCQ {//destripe_isk[7:4], 
                                          destripe_isk_q[0],
                                          destripe_isk[3:1]};
                  gt_rx_valid    <= #TCQ ~destripe_invalid;
                  end

        7'b0000100: begin // TWO_BIT_SHIFT
                  gt_rx_data     <= #TCQ {//destripe[63:32],
                                          destripe_q[15:0], 
                                          destripe[31:16]};
                  gt_rx_charisk  <= #TCQ {//destripe_isk[7:4],
                                          destripe_isk_q[1:0],
                                          destripe_isk[3:2]};
                  gt_rx_valid    <= #TCQ ~destripe_invalid;
                  end

        7'b0001000: begin // THREE_BIT_SHIFT
                        gt_rx_data     <= #TCQ {//destripe[63:32], 
                                                destripe_q[23:0],
                                                destripe[31:24]};
                        gt_rx_charisk  <= #TCQ {//destripe_isk[7:4], 
                                                destripe_isk_q[2:0],
                                                destripe_isk[3]};
                        gt_rx_valid    <= #TCQ ~destripe_invalid;
                        end
        
        7'b0010000: begin // pad bit insertion
                        gt_rx_data     <= #TCQ {//destripe[63:32], 
                                                pad[31:0]};
                        gt_rx_charisk  <= #TCQ {//destripe_isk[7:4], 
                                                pad_isk[3:0]};
                        gt_rx_valid    <= #TCQ ~destripe_invalid;
                        end

        default: begin
                 gt_rx_data     <= #TCQ destripe;
                 gt_rx_charisk  <= #TCQ destripe_isk;
                 gt_rx_valid    <= #TCQ ~destripe_invalid;
                 end

        endcase
      end else if ((LINK_WIDTH == 4)|| ((LINK_WIDTH == 2)&& !PPR_idle2_selected)) begin
        case (byte_alignment_nx_d)
        // If the alignngment is 4'b1000, then its possible there is another valid alignment
        // detected on this cycle
        4'b1000: begin
          gt_rx_data     <= #TCQ (multiple_alignments) ? {destripe[32+:32], pad} :
                                 (shift_align_b2b_cs)  ? {realign_bytes, destripe[0+:32]} :
                                                         destripe;
          gt_rx_charisk  <= #TCQ (multiple_alignments) ? {destripe_isk[4+:4], pad_isk} :
                                 (shift_align_b2b_cs)  ? {realign_isk, destripe_isk[0+:4]} :
                                                         destripe_isk;
          gt_rx_valid    <= #TCQ (multiple_alignments) ? {~destripe_invalid[4+:4], 4'b1111} :
                                 (shift_align_b2b_cs)  ? {realign_invalid, destripe_invalid[0+:4]} :
                                                          ~destripe_invalid;

          //*COVERAGE*
          //(cp_multiple_algins_8): See multiple alignments when the current alignment is 8
          //*COVERAGE*
          //(cp_shift_align_b2b_cs_8): See a back to back control symbol shift moving to alignment 8
          // only valid is 2 -> 8 based on striping requirements and cs lengths
        end
        // If the alignngment is 4'b0100, then its possible there is another valid alignment
        // detected on this cycle
        //FIXME
        4'b0100: begin
          gt_rx_data    <= #TCQ {realign_bytes[0+:24], destripe[24+:DATA_WIDTH-24]};
          gt_rx_charisk <= #TCQ {realign_isk[0+:3], destripe_isk[3+:CHARIS_WIDTH-3]};
          gt_rx_valid   <= #TCQ {~realign_invalid[0+:3], ~destripe_invalid[3+:CHARIS_WIDTH-3]};
          //*COVERAGE*
          //(cp_multiple_algins_4): See multiple alignments when the current alignment is 4
          //*COVERAGE*
          //(cp_shift_align_b2b_cs_4): See a back to back control symbol shift moving to alignment 4
          // only valid is 1 -> 4 based on striping requirements and cs lengths
        end
        4'b0010: begin
          gt_rx_data    <= #TCQ {realign_bytes[0+:16], destripe[16+:DATA_WIDTH-16]};
          gt_rx_charisk <= #TCQ {realign_isk[0+:2], destripe_isk[2+:CHARIS_WIDTH-2]};
          gt_rx_valid   <= #TCQ {~realign_invalid[0+:2], ~destripe_invalid[2+:CHARIS_WIDTH-2]};

        end
        4'b0001: begin
          gt_rx_data    <= #TCQ {realign_bytes[0+:8], destripe[8+:DATA_WIDTH-8]};
          gt_rx_charisk <= #TCQ {realign_isk[0+:1], destripe_isk[1+:CHARIS_WIDTH-1]};
          gt_rx_valid   <= #TCQ {~realign_invalid[0+:1], ~destripe_invalid[1+:CHARIS_WIDTH-1]};
        end
        default: begin
          gt_rx_data    <= #TCQ {DATA_WIDTH{1'bX}};
          gt_rx_charisk <= #TCQ {CHARIS_WIDTH{1'bX}};
          gt_rx_valid   <= #TCQ {CHARIS_WIDTH{1'bX}};
        end
        endcase
      end else if ((LINK_WIDTH == 2)&& PPR_idle2_selected) begin
        case (byte_alignment_2x_d) 
        11'b00000000001: begin // pass as is
                   gt_rx_data     <= #TCQ destripe;
                   gt_rx_charisk  <= #TCQ destripe_isk;
                   gt_rx_valid    <= #TCQ ~destripe_invalid;
                 end

        11'b00000000010: begin // strip last 2 bytes
                   gt_rx_data     <= #TCQ {destripe[63:16], pad[15:0]};
                   gt_rx_charisk  <= #TCQ {destripe_isk[7:2],pad_isk[1:0]};
                   gt_rx_valid    <= #TCQ ~destripe_invalid;
                 end

        11'b00000000100: begin // state s2
                   gt_rx_data     <= #TCQ {destripe[63:48], pad[15:0], destripe[47:16] };
                   gt_rx_charisk  <= #TCQ {destripe_isk[7:6],pad_isk[1:0], destripe_isk[5:2]};
                   gt_rx_valid    <= #TCQ ~destripe_invalid;
                 end

        11'b00000001000: begin // state s1
                   gt_rx_data     <= #TCQ {destripe_q[15:0], destripe[63:16]};
                   gt_rx_charisk  <= #TCQ {destripe_isk_q[1:0], destripe_isk[7:2]};
                   gt_rx_valid    <= #TCQ ~destripe_invalid;
                 end

        11'b00000010000: begin // state s3, condition 1, shifting from s2 to s3
                   gt_rx_data     <= #TCQ {destripe_q[15:0], destripe[63:16]};
                   gt_rx_charisk  <= #TCQ {destripe_isk_q[1:0], destripe_isk[7:2]};
                   gt_rx_valid    <= #TCQ ~destripe_invalid;
                 end

        11'b00000100000: begin // state s3, condition 2
                   gt_rx_data     <= #TCQ {destripe_q[15:0], destripe[63:48], destripe[31:0]};
                   gt_rx_charisk  <= #TCQ {destripe_isk_q[1:0], destripe_isk[7:6], destripe_isk[3:0]};
                   gt_rx_valid    <= #TCQ ~destripe_invalid;
                 end

        11'b00001000000: begin // state s3, transition to s1
                   gt_rx_data     <= #TCQ {destripe_q[15:0], destripe[63:16]};
                   gt_rx_charisk  <= #TCQ {destripe_isk_q[1:0], destripe_isk[7:2]};
                   gt_rx_valid    <= #TCQ ~destripe_invalid;
                 end

        11'b00010000000: begin // state s2, transition to ALIGN
                   gt_rx_data     <= #TCQ {destripe_q[15:0], destripe[63:48], destripe[31:0]};
                   gt_rx_charisk  <= #TCQ {destripe_isk_q[1:0], destripe_isk[7:6], destripe_isk[3:0]};
                   gt_rx_valid    <= #TCQ ~destripe_invalid;
                 end

        11'b00100000000: begin // state s2, transition to s0
                   gt_rx_data     <= #TCQ {destripe_q[15:0], destripe[63:48], destripe[31:0]};
                   gt_rx_charisk  <= #TCQ {destripe_isk_q[1:0], destripe_isk[7:6], destripe_isk[3:0]};
                   gt_rx_valid    <= #TCQ ~destripe_invalid;
                 end

        11'b01000000000: begin // state s2, transition to s1
                   gt_rx_data     <= #TCQ {destripe_q[15:0], destripe[63:16]};
                   gt_rx_charisk  <= #TCQ {destripe_isk_q[1:0], destripe_isk[7:2]};
                   gt_rx_valid    <= #TCQ ~destripe_invalid;
                 end

        default: begin
                 gt_rx_data     <= #TCQ destripe;
                 gt_rx_charisk  <= #TCQ destripe_isk;
                 gt_rx_valid    <= #TCQ ~destripe_invalid;
                 end

        endcase
      end
    end
  end

  //*COVERPOINT*
  //(cp_align_switch_x1_pre_init): cover that alignment switches for a x1 core before
  // port init.

  //*COVERPOINT*
  //(cp_align_switch_x2_pre_init): cover that alignment switches for a x2 core before
  // port init.

  //*COVERPOINT*
  //(cp_align_switch_x1_post_init): cover that alignment switches for a x1 core after
  // port init.

  //*COVERPOINT*
  //(cp_align_switch_x2_post_init): cover that alignment switches for a x2 core after
  // port init.
  // }}} Byte Alignment -------------------------

  // {{{ Clock Domain Crossing ------------------
  // For a x1 or x2 core, 4 and 8 bytes are received per cycles which can be directly shifted into 
  // a 64 bit data bus 
  generate if (LINK_WIDTH == 1 || LINK_WIDTH == 2) begin: ppr_out_x12_gen
    reg phy_rise_edge_det;
    reg phy_rise_edge_det_q;

    // Detect the rising edge of the phy clock
    always @(posedge phy_clk) begin
      if (phy_rst_q) begin
        phy_rise_edge_det <= #TCQ 1'b0;
      end else begin
        phy_rise_edge_det <= #TCQ ~phy_rise_edge_det;
      end
    end

    //Start out with 1 so the byte_idx will immediately load after a reset
    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        phy_rise_edge_det_q  <= #TCQ 1'b1;
      end else begin
        phy_rise_edge_det_q  <= #TCQ phy_rise_edge_det;
      end
    end

    wire phy_clk_edge_detected = phy_rise_edge_det_q != phy_rise_edge_det;

    // No reset needed since its not control
    always @(posedge gt_pcs_clk) begin
      if (phy_rst_q) begin            //9/24/2014, CR 824966, added default reset condition for below signals. 
        gt_rx_data_nx_q     <= #TCQ 0;//this is to make sure that at reset these signals are in known state.
        gt_rx_charisk_nx_q  <= #TCQ 0;
        gt_rx_valid_nx_q    <= #TCQ 0;
      end else if (PPI_mode_1x) begin
        gt_rx_data_nx_q     <= #TCQ {gt_rx_data_nx_q[31:0], gt_rx_data[31:0]};
        gt_rx_charisk_nx_q  <= #TCQ {gt_rx_charisk_nx_q[3:0], gt_rx_charisk[3:0]};
        gt_rx_valid_nx_q    <= #TCQ {gt_rx_valid_nx_q, &gt_rx_valid[3:0]};
      end else begin
        gt_rx_data_nx_q     <= #TCQ {gt_rx_data_nx_q, gt_rx_data};
        gt_rx_charisk_nx_q  <= #TCQ {gt_rx_charisk_nx_q, gt_rx_charisk};
        gt_rx_valid_nx_q    <= #TCQ {gt_rx_valid_nx_q, &gt_rx_valid};
      end
    end

  // For a x4 link width, 128 bits arrive at a time, so we need to only select
  // out 64 per phy clock cycle
  end else if (LINK_WIDTH == 4) begin: ppr_out_x4_gen
    reg gt_rise_edge_det;
    reg gt_rise_edge_det_q;

    // Detect the rising edge of the phy clock
    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        gt_rise_edge_det <= #TCQ 1'b0;
      end else begin
        gt_rise_edge_det <= #TCQ ~gt_rise_edge_det;
      end
    end

    //Start out with 1 so the byte_idx will immediately load after a reset
    always @(posedge phy_clk) begin
      if (phy_rst_q) begin
        gt_rise_edge_det_q  <= #TCQ 1'b1;
      end else begin
        gt_rise_edge_det_q  <= #TCQ gt_rise_edge_det;
      end
    end

    wire gt_clk_edge_detected = gt_rise_edge_det_q != gt_rise_edge_det;

    // Based on the link width increment through the byte locations
    // of the data in the phy clock domain. This is only needed for x1
    // cores where the gt_pcs_clk is faster than phy_clk. Because the edge 
    // detector will not be able to detect the rising edge until a cycle later, 
    // the load value of the byte counter will need to start at the second 
    // half of the dword.
    reg byte_idx;

    always @(posedge phy_clk) begin
      if (gt_clk_edge_detected) begin
        byte_idx <= #TCQ 0;
      end else begin
        byte_idx <= #TCQ 1;
      end
    end

    // Traindown register case
    always @(posedge gt_pcs_clk) begin
      if (gt_pcs_rst_q) begin
        gt_rx_valid_q       <= #TCQ 0;
        gt_rx_valid_1x_q    <= #TCQ 0;
      end else begin
        gt_rx_data_q        <= #TCQ gt_rx_data[31:0];
        gt_rx_charisk_q     <= #TCQ gt_rx_charisk[3:0];
        gt_rx_valid_q       <= #TCQ gt_rx_valid[3:0];

        gt_rx_data_1x_q     <= #TCQ {gt_rx_data_q[31:0], gt_rx_data[31:0]};
        gt_rx_charisk_1x_q  <= #TCQ {gt_rx_charisk_q[3:0], gt_rx_charisk[3:0]};
        gt_rx_valid_1x_q    <= #TCQ {&gt_rx_valid_q[3:0], &gt_rx_valid[3:0]};
      end
    end

    always @(posedge phy_clk) begin
      if (gt_pcs_rst_q) begin
        gt_rx_valid_nx_q    <= #TCQ 0;
      end else begin
        gt_rx_data_nx_q       <= #TCQ gt_rx_data[byte_idx*64+:64];
        gt_rx_charisk_nx_q    <= #TCQ gt_rx_charisk[byte_idx*8+:8];
        gt_rx_valid_nx_q      <= #TCQ gt_rx_valid[byte_idx*2+:2];
      end
    end
  end endgenerate

  // Register the data in the PHY clock domain
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PPR_rx_data         <= #TCQ 0;
      PPR_rx_charisk      <= #TCQ 0;
      PPR_rx_valid        <= #TCQ 0;
      PPR_out_of_sync     <= #TCQ 1;
    end else begin
      // Train down case for x4
      if (PPI_mode_1x && LINK_WIDTH == 4) begin
        PPR_rx_data         <= #TCQ {PPR_rx_data, gt_rx_data_1x_q};
        PPR_rx_charisk      <= #TCQ {PPR_rx_charisk, gt_rx_charisk_1x_q};
        PPR_rx_valid        <= #TCQ {PPR_rx_valid, gt_rx_valid_1x_q};
        PPR_out_of_sync     <= #TCQ gt_out_of_sync;
 
      // Train down case for x2
      end else if (PPI_mode_1x && LINK_WIDTH == 2) begin
        PPR_rx_data         <= #TCQ {PPR_rx_data, gt_rx_data_nx_q};
        PPR_rx_charisk      <= #TCQ {PPR_rx_charisk, gt_rx_charisk_nx_q};
        PPR_rx_valid        <= #TCQ {PPR_rx_valid, gt_rx_valid_nx_q};
        PPR_out_of_sync     <= #TCQ gt_out_of_sync;

      end else begin
        PPR_rx_data         <= #TCQ gt_rx_data_nx_q;
        PPR_rx_charisk      <= #TCQ gt_rx_charisk_nx_q;
        PPR_rx_valid        <= #TCQ gt_rx_valid_nx_q;
        PPR_out_of_sync     <= #TCQ gt_out_of_sync;
      end
    end
  end
  // }}} end Clock Domain Crossing

//_________
  //State Machine States
  localparam ALIGN = 3'd0;
  localparam S0    = 3'd1;
  localparam S1    = 3'd2;
  localparam S2    = 3'd3;
  localparam S3    = 3'd4;
//______________________________________________________________________________

  
//______________________________________________________________________________

    `ifdef SIMULATION
    reg [20*8-1:0] rx_align_next_state_string = "null";
    reg [20*8-1:0] rx_align_state_string      = "null";

    always @* begin
      case (rx_align_state)
        ALIGN:          rx_align_state_string = "ALIGN";
        S0:             rx_align_state_string = "S0";
        S1:             rx_align_state_string = "S1";
        S2:             rx_align_state_string = "S2";
        S3:             rx_align_state_string = "S3";
        default:        rx_align_state_string = "INVALID";
      endcase
      case (rx_align_next_state)
        ALIGN:          rx_align_next_state_string = "ALIGN";
        S0:             rx_align_next_state_string = "S0";
        S1:             rx_align_next_state_string = "S1";
        S2:             rx_align_next_state_string = "S2";
        S3:             rx_align_next_state_string = "S3";
        default:        rx_align_next_state_string = "INVALID";
      endcase
    end
  `endif
//______________________________________________________________________________
wire [2:0] destripe_pdsc_add;
wire sop_hunt_2x;
reg  [2:0] destripe_pdsc_add_reg; 
wire bit_7;
wire bit_5;
wire bit_3;
wire bit_1;
wire bit_11;
wire bit_31;
wire bit_51;
wire bit_71;
reg  bit_lsb_lw_misalign; 
reg  bit_lsb_lw_align   ; 
reg  bit_msb_up_misalign; 
reg  bit_msb_up_align   ; 

assign destripe_pdsc_add[0] = destripe_pdsc[7] ||
                              destripe_pdsc[5] ||
                              destripe_pdsc[3] ||
                              destripe_pdsc[1];

  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) 
      destripe_pdsc_add_reg <= #TCQ 3'b0;
    else if (!PPI_port_initialized)
      destripe_pdsc_add_reg <= #TCQ 3'b0;
    else 
      destripe_pdsc_add_reg <= #TCQ destripe_pdsc_add;
  end

  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      csymbol_monitor_2x <= #TCQ 1;
    end else begin
      if (!PPI_port_initialized) begin
        csymbol_monitor_2x <= #TCQ 1;
      end else if (LINK_WIDTH == 2) begin
        if (|destripe_pdsc && csymbol_monitor_2x) begin
          csymbol_monitor_2x <= #TCQ 0;
        end
    end
  end
  end
// check for SOP for new packet
assign sop_hunt_2x = csymbol_monitor_2x || destripe_pdsc_add[0] || bit_msb_up_align;


    always @(destripe_pdsc) begin
      casex ({destripe_pdsc[7], 
             destripe_pdsc[5],
             destripe_pdsc[3],
             destripe_pdsc[1]})
        4'bxxx1: begin
                 bit_lsb_lw_misalign = 1'b1;
                 bit_lsb_lw_align    = 1'b0;
                 bit_msb_up_misalign = 1'b0;
                 bit_msb_up_align    = 1'b0;
                 end
        4'bxx10: begin
                 bit_lsb_lw_misalign = 1'b0;
                 bit_lsb_lw_align    = 1'b1;
                 bit_msb_up_misalign = 1'b0;
                 bit_msb_up_align    = 1'b0;
                 end
        4'bx100: begin
                 bit_lsb_lw_misalign = 1'b0;
                 bit_lsb_lw_align    = 1'b0;
                 bit_msb_up_misalign = 1'b1;
                 bit_msb_up_align    = 1'b0;
                 end
        4'b1000: begin
                 bit_lsb_lw_misalign = 1'b0;
                 bit_lsb_lw_align    = 1'b0;
                 bit_msb_up_misalign = 1'b0;
                 bit_msb_up_align    = 1'b1;
                 end
        default: begin
                 bit_lsb_lw_misalign = 1'b0;
                 bit_lsb_lw_align    = 1'b0;
                 bit_msb_up_misalign = 1'b0;
                 bit_msb_up_align    = 1'b0;
                 end
      endcase
    end

assign bit_11 = bit_lsb_lw_misalign && sop_hunt_2x && !csymbol_monitor_2x;
assign bit_31 = bit_lsb_lw_align    && sop_hunt_2x && !csymbol_monitor_2x;   
assign bit_51 = bit_msb_up_misalign && sop_hunt_2x && !csymbol_monitor_2x;
assign bit_71 = bit_msb_up_align    && sop_hunt_2x && !csymbol_monitor_2x;   


assign bit_7 = (sop_hunt_2x && csymbol_monitor_2x && destripe_pdsc[7])
               || bit_71;
assign bit_5 = (sop_hunt_2x && csymbol_monitor_2x && destripe_pdsc[5])
               || bit_51;
assign bit_3 = (sop_hunt_2x && csymbol_monitor_2x && destripe_pdsc[3])
               || bit_31;
assign bit_1 = (sop_hunt_2x && csymbol_monitor_2x && destripe_pdsc[1])
               || bit_11;

//______________________________________________________________________________
  always @(posedge gt_pcs_clk)
  begin
    if (gt_pcs_rst_q)
        begin
          rx_align_state <= #TCQ ALIGN;
        end
    else
        begin
          rx_align_state <= #TCQ rx_align_next_state;
        end
  end
//______________________________________________________________________________
  always @(*)
  begin
    //Set Initial defaults
    byte_alignment_2x_d = 11'b00000000001;

    case (rx_align_state)
       ALIGN:begin
                if (bit_5) begin
                  rx_align_next_state = S2;                   // 6th bit is PDSC
                  byte_alignment_2x_d = 11'b00000000100;
                  end
                else if (bit_1) begin
                  rx_align_next_state = S0;                   // 2nd bit is PDSC
                  byte_alignment_2x_d = 11'b00000000010;
                  end
                else begin
                  rx_align_next_state = ALIGN;                // align state only
                  byte_alignment_2x_d = 11'b00000000001;
                end
             end

       S0:begin // 2nd bit is PDSC
                  rx_align_next_state = S1;                   // 2nd bit is PDSC
                  byte_alignment_2x_d = 11'b00000001000;
            end

       S1:begin // 2nd bit is PDSC
                if (bit_7 || bit_3) begin
                  rx_align_next_state = ALIGN;                // 7th, 1st bit is PDSC
                  byte_alignment_2x_d = 11'b00000000001;
                  end
                else if (bit_5) begin
                  rx_align_next_state = S3;                   // 6th bit is PDSC
                  byte_alignment_2x_d = 11'b00000010000;
                  end
                else begin
                  rx_align_next_state = S1;                   // 2nd bit is PDSC
                  byte_alignment_2x_d = 11'b00000001000;
                end
            end

       S2:begin // 6th bit is PDSC
                if (bit_3) begin
                  rx_align_next_state = ALIGN;            
                  byte_alignment_2x_d = 11'b00010000000;
                  end 
                else if (bit_1) begin
                  rx_align_next_state = S1;
                  byte_alignment_2x_d = 11'b01000000000;
                end
                else begin
                  rx_align_next_state = S3;                   // 6th bit is PDSC
                  byte_alignment_2x_d = 11'b00000010000;
                end
            end

       S3:begin // 6th bit is PDSC
                if (bit_7 || bit_3) begin
                  rx_align_next_state = ALIGN;                // 7th, 1st bit is PDSC
                  if (bit_7)
                    byte_alignment_2x_d = 11'b00000000001;               
                  else if (bit_3)
                    byte_alignment_2x_d = 11'b00000100000;             
                end
                else if (bit_1) begin
                  rx_align_next_state = S1;                   // 2nd bit is PDSC
                  byte_alignment_2x_d = 11'b00001000000;
                end
                else begin
                  rx_align_next_state = S3;                   // 6th bit is PDSC
                  byte_alignment_2x_d = 11'b00000010000;
                end 
            end

       default: begin
                     byte_alignment_2x_d = 11'b00000000001;
		             rx_align_next_state = ALIGN; //7/20/2014, added to avoide latch
                end

   endcase
  end
//______________________________________________________________________________
//______________________________________________________________________________
 

    `ifdef SIMULATION
    reg [20*8-1:0] rx_1x_align_next_state_string = "null";
    reg [20*8-1:0] rx_1x_align_state_string      = "null";

    always @* begin
      case (rx_1x_align_state)
        ALIGN:             rx_1x_align_state_string = "ALIGN_1X";
        ONE_BIT_SHIFT:     rx_1x_align_state_string = "ONE_BIT_SHIFT";
        TWO_BIT_SHIFT:     rx_1x_align_state_string = "TWO_BIT_SHIFT";
        THREE_BIT_SHIFT:   rx_1x_align_state_string = "THREE_BIT_SHIFT";
        INTER_STATE:       rx_1x_align_state_string = "INTER_STATE";
        INTER_STATE2:       rx_1x_align_state_string = "INTER_STATE2";
        INTER_STATE1:       rx_1x_align_state_string = "INTER_STATE1";
        default:           rx_1x_align_state_string = "INVALID";
      endcase
      case (rx_1x_align_next_state)
        ALIGN:             rx_1x_align_next_state_string = "ALIGN_1X";
        ONE_BIT_SHIFT:     rx_1x_align_next_state_string = "ONE_BIT_SHIFT";
        TWO_BIT_SHIFT:     rx_1x_align_next_state_string = "TWO_BIT_SHIFT";
        THREE_BIT_SHIFT:   rx_1x_align_next_state_string = "THREE_BIT_SHIFT";
        INTER_STATE:       rx_1x_align_next_state_string = "INTER_STATE";
        INTER_STATE2:       rx_1x_align_next_state_string = "INTER_STATE2";
        INTER_STATE1:       rx_1x_align_next_state_string = "INTER_STATE1";
        default:           rx_1x_align_next_state_string = "INVALID";
      endcase
    end
  `endif

//____ below code is for 1x mode _______________________________________________

reg bit_3_1x;
reg bit_2_1x;
reg bit_1_1x;
reg bit_0_1x;
// below mux logic is to find SOP of next packet
    always @(destripe_pdsc) begin // this code looks for SOP from lower to upper bits
      casex ({destripe_pdsc[3], 
              destripe_pdsc[2],
              destripe_pdsc[1],
              destripe_pdsc[0]})

	     4'bxxx1: begin 
                     bit_3_1x = 1'b0;
                     bit_2_1x = 1'b0;
                     bit_1_1x = 1'b0;
                     bit_0_1x = 1'b1;
             end

	     4'bxx10: begin 
                     bit_3_1x = 1'b0;
                     bit_2_1x = 1'b0;
                     bit_1_1x = 1'b1;
                     bit_0_1x = 1'b0;
             end

	     4'bx100: begin 
                     bit_3_1x = 1'b0;
                     bit_2_1x = 1'b1;
                     bit_1_1x = 1'b0;
                     bit_0_1x = 1'b0;
             end

	     4'b1000: begin 
                     bit_3_1x = 1'b1;
                     bit_2_1x = 1'b0;
                     bit_1_1x = 1'b0;
                     bit_0_1x = 1'b0;
             end
             
             default: begin
                     bit_3_1x = 1'b0;
                     bit_2_1x = 1'b0;
                     bit_1_1x = 1'b0;
                     bit_0_1x = 1'b0;
             end
         endcase
      end

// logic to get the  csymbol_monitor_1x
  always @(posedge gt_pcs_clk) begin
    if (gt_pcs_rst_q) begin
      csymbol_monitor_1x <= #TCQ 1;
    end else begin
      if (!PPI_port_initialized) begin
        csymbol_monitor_1x <= #TCQ 1;
      end else if (LINK_WIDTH == 1 || PPI_mode_1x) begin
        if (|destripe_pdsc && csymbol_monitor_1x) begin
          csymbol_monitor_1x <= #TCQ 0;
        end
    end
  end
  end

wire sop_hunt_1x;
reg sop_hunt_1x_q;
wire [2:0] add_lower_nibble;
reg  [2:0] add_lower_nibble_q;
reg bit_3_1x_q;
reg bit_2_1x_q;
reg bit_1_1x_q;
reg bit_0_1x_q;
reg bit_2_1x_q1;
reg bit_1_1x_q1 ;
reg sync_1x_q;
reg sync_latch;
reg reset_sync_latch;
reg sync_latch_q;
reg sync_latch_q1;
wire sync_1x;
wire sync_det;

always @(posedge gt_pcs_clk) begin
  if (gt_pcs_rst_q) begin
    bit_3_1x_q <= #TCQ 0 ;
    bit_2_1x_q <= #TCQ 0 ; 
    bit_1_1x_q <= #TCQ 0 ;
    bit_0_1x_q <= #TCQ 0 ;
    bit_2_1x_q1 <= #TCQ 0 ;
    bit_1_1x_q1 <= #TCQ 0 ;
    sync_latch_q <= #TCQ 0;
    sync_latch_q1 <= #TCQ 0;
  end else begin
    bit_3_1x_q <= #TCQ bit_3_1x;
    bit_2_1x_q <= #TCQ bit_2_1x;
    bit_1_1x_q <= #TCQ bit_1_1x;
    bit_2_1x_q1 <= #TCQ bit_2_1x_q;
    bit_1_1x_q1 <= #TCQ bit_1_1x_q;
    bit_0_1x_q <= #TCQ bit_0_1x;
    sync_latch_q <= #TCQ sync_latch;
    sync_latch_q1 <= #TCQ sync_latch_q;
  end
end

//______________________________________________________________________________

//______________________________________________________________________________

assign sync_det = (    (destripe_isk[3] && destripe[31:24]==8'h3c)
            || (destripe_isk[2] && destripe[23:16]==8'h3c)
	    || (destripe_isk[1] && destripe[15:8] ==8'h3c)
	    || (destripe_isk[0] && destripe[7:0]  ==8'h3c)
	  );

always @(posedge gt_pcs_clk)
begin
  if (gt_pcs_rst_q)
      begin
        add_lower_nibble_q <= #TCQ 3'b0;   
      end
  else if ( sync_det === 1'b1 && sop_hunt_1x_q == 1'b0) 
      begin
        add_lower_nibble_q <= #TCQ 3'b0;   
      end
  else
      begin
        add_lower_nibble_q <= #TCQ add_lower_nibble;   
      end
end

assign add_lower_nibble = (destripe_pdsc[3] +
                           destripe_pdsc[2] +
                           destripe_pdsc[1] +
                           destripe_pdsc[0] +
                           (add_lower_nibble_q[0] && PPR_idle2_selected)
                            );


assign sop_hunt_1x = !PPI_port_initialized ? 1'b1 :
                                          //sop_hunt_1x_q ? 1'b0 :
                                          (add_lower_nibble[0]);

always @(posedge gt_pcs_clk) begin
  if (gt_pcs_rst_q) begin
    sop_hunt_1x_q <= #TCQ 0;
  end else begin
    sop_hunt_1x_q <= #TCQ sync_det;
  end
end



wire bit_33_1x;
wire bit_22_1x;
wire bit_11_1x;
wire bit_00_1x;

assign bit_33_1x = bit_3_1x && sop_hunt_1x; // this is to test every new SOP
assign bit_22_1x = bit_2_1x && sop_hunt_1x; // -- " --
assign bit_11_1x = bit_1_1x && sop_hunt_1x; // -- " --
assign bit_00_1x = bit_0_1x && sop_hunt_1x; // -- " -- 

//___________________1x present state to next state converter __________________

  always @(posedge gt_pcs_clk)
  begin
    if (gt_pcs_rst_q)
        begin
          rx_1x_align_state <= #TCQ ALIGN_1X;
        end
    else
        begin
          rx_1x_align_state <= #TCQ rx_1x_align_next_state;
        end
  end

//________________Rx 1x state machine __________________________________________
  always @(*)
  begin
    case (rx_1x_align_state)
              ALIGN_1X: begin // no need to check any existing pdsc's
			                  if (bit_22_1x) begin            //0100
                                  rx_1x_align_next_state = THREE_BIT_SHIFT;
                                  byte_alignment_1x_d = 7'b0010000;
                              end else if (bit_11_1x) begin   //0010
                                  rx_1x_align_next_state = TWO_BIT_SHIFT;
                                  byte_alignment_1x_d = 7'b0010000;
                              end else if (bit_00_1x) begin    //0001
                                  rx_1x_align_next_state = ONE_BIT_SHIFT;
                                  byte_alignment_1x_d = 7'b0010000;
                              end else begin                   //1000
                                 rx_1x_align_next_state = ALIGN_1X;
                                 byte_alignment_1x_d = 7'b0000001;
                              end
                        end

       THREE_BIT_SHIFT: begin
      			            if (bit_33_1x) begin                                // completed earlier one 
                                    rx_1x_align_next_state = ALIGN_1X;          // and looking for fresh one
                                    byte_alignment_1x_d = 7'b0000001;
                            end else if (bit_11_1x && !destripe_pdsc[3]) begin  // completed earlier one    
                                    rx_1x_align_next_state = TWO_BIT_SHIFT;     // and looking for fresh one
                                    byte_alignment_1x_d = 7'b0010000;
                            end else if (bit_00_1x && !destripe_pdsc[3]) begin  // completed earlier one    
                                    rx_1x_align_next_state = ONE_BIT_SHIFT;     // and looking for fresh one
                                    byte_alignment_1x_d = 7'b0010000;
                            end else if (bit_11_1x && destripe_pdsc[3]) begin   // first one is present    
                                    rx_1x_align_next_state = INTER_STATE;       // and 2nd transaction came
                                    byte_alignment_1x_d = 7'b0001000;             // but no pure back to back
                            end else if (bit_00_1x && destripe_pdsc[3]) begin   // first one is present    
                                    rx_1x_align_next_state = INTER_STATE;       // and 2nd transaction came
                                    byte_alignment_1x_d    = 7'b0001000;
                            end else begin
                                    rx_1x_align_next_state = THREE_BIT_SHIFT;
                                    byte_alignment_1x_d = 7'b0001000;
                            end
                     end

       TWO_BIT_SHIFT: begin 
			                  if (bit_33_1x) begin // fresh transaction
                                      rx_1x_align_next_state = ALIGN_1X;
                                      byte_alignment_1x_d = 7'b0000001;
                              end else if (bit_22_1x) begin // fresh transaction
                                      rx_1x_align_next_state = THREE_BIT_SHIFT;
                                      byte_alignment_1x_d = 7'b0010000;
                              end else if (bit_00_1x && !destripe_pdsc[2]) begin // fresh transaction
                                      rx_1x_align_next_state = ONE_BIT_SHIFT;
                                      byte_alignment_1x_d = 7'b0010000;
                              end else if (bit_00_1x && destripe_pdsc[2]) begin
                                      rx_1x_align_next_state = INTER_STATE2;
                                      byte_alignment_1x_d    = 7'b0000100;
                              end else begin
                                      rx_1x_align_next_state = TWO_BIT_SHIFT;
                                      byte_alignment_1x_d = 7'b0000100;
                              end
                     end

       ONE_BIT_SHIFT: begin 
			                if (bit_33_1x) begin
                                    rx_1x_align_next_state = ALIGN_1X;
                                    byte_alignment_1x_d = 7'b0000001;
                            end else if (bit_22_1x) begin
                                    rx_1x_align_next_state = THREE_BIT_SHIFT;
                                    byte_alignment_1x_d = 7'b0010000;
                            end else if (bit_11_1x) begin
                                    rx_1x_align_next_state = TWO_BIT_SHIFT;
                                    byte_alignment_1x_d = 7'b0010000;
                            end else begin
                                    rx_1x_align_next_state = ONE_BIT_SHIFT;
                                    byte_alignment_1x_d = 7'b0000010;
                            end
                      end


       INTER_STATE: begin
                        if (destripe_pdsc_q[1]) begin          // this is for 2 bit shift
                                rx_1x_align_next_state = TWO_BIT_SHIFT;
                                byte_alignment_1x_d = 7'b0000100;
                        end else if (destripe_pdsc_q[0]) begin // this is for 1 bit shift
                                rx_1x_align_next_state = ONE_BIT_SHIFT;
                                byte_alignment_1x_d = 7'b0000010;
                        end else begin // below updates to remove latch
 			                    rx_1x_align_next_state = ALIGN_1X;//7/20/2014
			                    byte_alignment_1x_d = 7'b0000001;//7/20/2014
                        end
                    end

       INTER_STATE2: begin
                          rx_1x_align_next_state = ONE_BIT_SHIFT;
                          byte_alignment_1x_d = 7'b0000010;
                     end

       default: begin
                     rx_1x_align_next_state = ALIGN_1X;
                     byte_alignment_1x_d    = 7'b0000001;
                end
    endcase
  end
//______________________________________________________________________________

endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//---------------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/phy/srio_gen2_v4_1_16_phy_top.v#1 $
//---------------------------------------------------------------------------
`timescale 1ps/1ps
// ------------------------------------------------
// below attribute is added to supress the synthesis warnings in vivado tool 8:3332
(* DowngradeIPIdentifiedWarnings="yes" *)
// ------------------------------------------------


module srio_gen2_v4_1_16_phy_top
#(parameter TCQ           = 100,        // in ps
  parameter SIM_TRAIN     = 0,          // Allows fast train {0:FULL, 1:FAST, 2:TRAINED}
  parameter LINK_WIDTH    = 1,          // Number of GT lanes {1, 2, 4}
  parameter MODE_XG       = 5,          // Line rates {1/1.25, 2/2.5, 3/3.125, 5/5, 6/6.25}
  parameter IDLE1         = 1,          // Include the IDLE1 sequence {0,1}
  parameter IDLE2         = 0,          // Include the IDLE2 sequence {0,1}
  parameter SCRAM         = 0,          // Inserts the scrambler modules {0,1}
  parameter VC            = 0,          // Highest number VC supported {0,1}
  parameter RETRY         = 1,          // Includes Retry protocol {0, 1}
  parameter LINK_REQUESTS = 3,          // Additional link requests to send prior to port_error {0-6,7/inf}
  parameter TARGET_DS     = 0,          // Additional link requests to send prior to port_error {0-6,7/inf}
  parameter PHY_EF_PTR    = 16'h0100,   // Location of PHY  ext features {0x100+}
  parameter LANE_EF_PTR   = 16'h0400,   // Location of Lane ext features {0x400+}
  parameter VC_EF_PTR     = 16'h0800,   // Location of VC   ext features {0x800+} (only if VC==1)
  parameter LINK_TIMEOUT  = 24'hFF_FFFF,// Link timeout ctr {0x000000-0xffffff}
  parameter PORT_TIMEOUT  = 24'hFF_FFFF,// Port timeout ctr {0x000000-0xffffff}
  parameter IS_HOST       = 1,          // Default Host value {0,1}
  parameter MASTER_EN     = 1,          // Default Master enable value {0,1}
  parameter DISCOVERED    = 0,          // Default discovered value {0,1}
  parameter DEBUG         = 0,          // Default discovered value {0,1}
  parameter VC1_CT        = 1,          // Default traffic mode for VC1 {0,1/continous}
  parameter USER_EF_PTR   = 16'h0000,   // Location of User ext features {0x0000 or 0x0900+}
  parameter SW_CSR        = 0,          // SW assisted error recovery enabled {0,1}
  parameter EVAL          = 1,          // Indicates an Evaluation Core
  parameter SWITCH_MODE   = 0,          // If the core is generated with Switch Mode Support
  parameter GT_BYTES      = 4           // Bytes on the GT Interface
)
 // {{{ ports -------------------------------------------------
 (input                              phy_clk,                    // PHY interface clock
  input                              phy_rst,                    // Reset for PHY clock Domain
  input                              log_clk,                    // LOG interface clock
  input                              log_rst,                    // Reset for LOG clock Domain
  input                              gt_pcs_clk,                 // GT Interface user clock
  input                              gt_pcs_rst,                 // Reset for GT clk domain
  input                              cfg_clk,                    // CFG Interface user clock
  input                              cfg_rst,                    // Reset for CFG clk domain
  input                              sim_train_en,               // Enable SIM_TRAIN mode for imp.
  input                              BT_phyt_tvalid,             // Valid data indicator
  output                             PT_phyt_tready,             // Destination Ready
  input  [63:0]                      BT_phyt_tdata,              // Packet for transfer
  input  [7:0]                       BT_phyt_tkeep,              // Byte Enable for transferred packet
  input                              BT_phyt_tlast,              // Last DW of incoming packet
  input  [7:0]                       BT_phyt_tuser,              // {1'b0, SKIP_CRC, 2'b00, VC, CRF, SRC_DSC}
  output [5:0]                       PT_phy_next_fm,             // Next packet's ackID
  output [5:0]                       PR_phy_last_ack,            // Last PA received by the PHY core
  input  [5:0]                       BR_phy_buf_stat,            // Buffer status from the RX buffer to be transmitted
  input                              UG_phy_mce,                 // Send MCE control symbol
  input                              UG_phy_link_reset,          // Send link reset control symbols
  output                             PR_link_initialized,        // Indicates we are ready to transmit data
  output                             PR_phyr_tvalid,             // Valid data indicator
  input                              BR_phyr_tready,             // Destination Ready
  output [63:0]                      PR_phyr_tdata,              // Packet for transfer
  output [7:0]                       PR_phyr_tkeep,              // Byte Enable for transferred packet
  output                             PR_phyr_tlast,              // Last DW of incoming packet
  output [7:0]                       PR_phyr_tuser,              // {5'h00, VC, CRF, src_dsc}
  output                             PT_phy_rewind,              // An error or retry condition is in progress
  output [5:0]                       PR_phy_rcvd_buf_stat,       // Buffer status received from the link partner
  output                             PR_phy_rcvd_mce,            // MCE control symbol received
  output                             PR_phy_rcvd_link_reset,     // Received 4 consecutive link reset control symbols
  output                             PR_port_error,              // Indicator that OLLM RX is in Port Error State
  output                             PP_port_initialized,        // Indicates port is initialized
  output                             PP_mode_1x,                 // Indicates the link trained down to 1x
  output                             PP_idle2_selected,          // Indicates the link is operating in IDLE2 mode
  output                             PP_idle_selected,           // Indicates the IDLE Sequence is selected
  input                              UG_force_reinit,            // Force reinitialization
  output [23:0]                      PC_port_timeout,            // Timeout value user can use to detect lost packet
  output                             PC_srio_host,               // Endpoint is the system host
  output                             PC_master_enable,           // Enable Request transactions
  input                              BT_tx_flow_control,         // Port negotiated to tx flow control
  output                             PC_maint_only,              // LOG can only send maintenance packets
  input                              CF_cfgp_awvalid,            // Write Command Valid
  output                             PC_cfgp_awready,            // Write Port Ready
  input  [23:0]                      CF_cfgp_awaddr,             // Write Address
  input                              CF_cfgp_wvalid,             // Write Data Valid
  output                             PC_cfgp_wready,             // Write Port Ready
  input  [31:0]                      CF_cfgp_wdata,              // Write Data
  input  [3:0]                       CF_cfgp_wstrb,              // Write Data byte enables
  output                             PC_cfgp_bvalid,             // Write Response Valid
  input                              CF_cfgp_bready,             // Write Response Fabric Ready
  input                              CF_cfgp_arvalid,            // Read Command Valid
  output                             PC_cfgp_arready,            // Read Port Ready
  input  [23:0]                      CF_cfgp_araddr,             // Read Address
  output                             PC_cfgp_rvalid,             // Read Response Valid
  input                              CF_cfgp_rready,             // Read Response Fabric Ready
  output [31:0]                      PC_cfgp_rdata,              // Read Data
  output [LINK_WIDTH*GT_BYTES*8-1:0] PP_gttx_data,               // Transmit Data to the GTs
  output [LINK_WIDTH*GT_BYTES-1:0]   PP_gttx_charisk,            // Transmit char is K to the GTs
  input  [LINK_WIDTH*GT_BYTES*8-1:0] GT_gtrx_data,               // Receive Data from the GTs
  input  [LINK_WIDTH*GT_BYTES-1:0]   GT_gtrx_charisk,            // Receive Data is K from the GTs
  input  [LINK_WIDTH*GT_BYTES-1:0]   GT_gtrx_chariscomma,        // Receive Data is comma
  input  [LINK_WIDTH*GT_BYTES-1:0]   GT_gtrx_disperr,            // Receive Data contains disperity Error
  input  [LINK_WIDTH*GT_BYTES-1:0]   GT_gtrx_notintable,         // Receive Data contains a not in table Error
  output [LINK_WIDTH-1:0]            PP_gttx_inhibit,            // TX Inhibit to the GTs
  input  [LINK_WIDTH-1:0]            GT_gtrx_chanisaligned,      // RX chanel is aligned across all GTs
  input                              GT_gtrx_reset_req,          // RX Buffer Error from the GTs
  input  [LINK_WIDTH-1:0]            GT_gtrx_reset_done,         // RX Buffer Reset Done
  output                             PP_gtrx_reset,              // Reset the GTs RX Buffer
  output                             PP_rx_lane_r,               // Receiving Data on lane R
  output                             PP_gtrx_chanbonden,         // Enable chanel bonding
  output [95:0]                      PP_debug,                   // Debugs from OPLM
  output [63:0]                      PT_debug,                   // Debugs from OLLM TX
  output [63:0]                      PR_debug                    // Debugs from OLLM RX
  );
  // }}} --------------------------------------------

  // {{{ Between the OPLM and OLLM_TX
  wire [63:0]                    PT_tx_data;
  wire [7:0]                     PT_tx_charisk;
  wire [1:0]                     PT_tx_valid;
  wire [1:0]                     PT_tx_early_valid;
  wire                           PT_tx_early_lreq;
  wire                           PP_ccomp_req;
  wire                           PT_ccomp_grant;
  wire                           PT_send_lreq;
  wire                           PP_lreq_sent;
  wire                           PP_out_of_sync;
  // }}}

  // {{{ Between the OPLM and the OLLM_RX
  wire [63:0]                    PP_rx_data;
  wire [7:0]                     PP_rx_charisk;
  wire [1:0]                     PP_rx_valid;
  // }}}

  // {{{ Between the OLLM_TX and OLLM_RX
  wire                           PT_sent_init_cs;
  wire                           PR_rewind;
  wire                           PR_send_rfr;
  wire                           PT_rfr_sent;

  wire                           PR_send_lreq;
  wire                           PR_send_pna;
  wire                           PT_lreq_sent;
  wire                           PT_pna_sent;
  wire                           PR_send_pr;
  wire                           PT_pr_sent;
  wire                           PR_send_lresp;
  wire                           PT_lresp_sent;
  wire [5:0]                     PR_last_good_pkt;
  wire [4:0]                     PR_cause;
  wire [4:0]                     PR_port_stat;
  wire                           PT_switch_crc_err;
  wire                           PR_rcvd_error_free_status;
  wire                           PT_sample_next_fm;
  // }}}

  // {{{ Between the OPLM and PHY_CFG
  wire                           PC_scram_disable;
  wire                           PC_force_1x;
  wire [2:0]                     PC_force_lane;
  wire                           PC_port_disable;
  wire                           PC_idle2_enable;
  wire [LINK_WIDTH*2-1:0]        PP_gtrx_tap_m1_status;
  wire [LINK_WIDTH*2-1:0]        PP_gtrx_tap_p1_status;
  wire [LINK_WIDTH-1:0]          PP_rx_scram_en;
  wire [LINK_WIDTH-1:0]          PP_receiver_trained;
  wire [LINK_WIDTH-1:0]          PP_idle2_rcvd;
  wire [LINK_WIDTH*4-1:0]        PP_rx_lane_number;
  wire [LINK_WIDTH*3-1:0]        PP_rx_port_width;
  wire [LINK_WIDTH*4-1:0]        PP_gt_decode_error;
  wire [LINK_WIDTH-1:0]          PP_lane_sync;
  // }}}

  // {{{ Between the OLLM_TX and PHY_CFG
  wire                           PC_send_lreq;
  wire [2:0]                     PC_lreq_cmd;
  wire [5:0]                     PC_next_fm;
  wire [4:0]                     PR_rcvd_port_stat;
  // }}} End ollm_tx_top signals

  // {{{ Between the OLLM_RX and PHY_CFG
  wire [5:0]                     PR_next_rcvd_pkt;
  wire [5:0]                     PC_next_rcvd_pkt;
  wire [5:0]                     PC_last_ack;
  wire                           PR_rcvd_lresp;
  wire [5:0]                     PR_ackid_status;
  wire [23:0]                    PC_link_timeout;
  wire                           PR_output_retry_stop;
  wire                           PR_output_error_stop;
  wire                           PR_input_retry_stop;
  wire                           PR_input_error_stop;
  wire                           PR_rcvd_pa_or_pna;
  wire                           PC_clr_port_error;
  wire                           PC_input_maint_only;
  wire                           PC_error_disable;
  wire                           PC_vc_ct;
  wire                           PC_load_nextpkt;
  // }}}

  // {{{ Between multiple blocks and the PHY_CFG
  wire                           PC_load_ackids;
  wire                           PC_vc_en;
  // }}}


  // {{{ Core stats assignment - can't find a better place for this
  wire  PHY_core_stats_info = {63'h0,
                                PR_send_pna};
  // }}}


  // {{{ oplm_top instantiation
  //--------------------------------------------
  srio_gen2_v4_1_16_oplm_top
    #(.TCQ                       (TCQ),
      .LINK_WIDTH                (LINK_WIDTH),
      .IDLE1                     (IDLE1),
      .IDLE2                     (IDLE2),
      .MODE_XG                   (MODE_XG),
      .SCRAM                     (SCRAM),
      .SIM_TRAIN                 (SIM_TRAIN),
      .GT_BYTES                  (GT_BYTES),
      .DEBUG                     (DEBUG),
      .EVAL                      (EVAL))
    oplm_top_inst
     (.gt_pcs_clk                (gt_pcs_clk),
      .gt_pcs_rst                (gt_pcs_rst),
      .phy_clk                   (phy_clk),
      .phy_rst                   (phy_rst),
      .sim_train_en              (sim_train_en),
      .UG_force_reinit           (UG_force_reinit),
      .PT_tx_data                (PT_tx_data),
      .PT_tx_charisk             (PT_tx_charisk),
      .PT_tx_valid               (PT_tx_valid),
      .PT_tx_early_lreq          (PT_tx_early_lreq),
      .PP_port_initialized       (PP_port_initialized),
      .PP_ccomp_req              (PP_ccomp_req),
      .PT_ccomp_grant            (PT_ccomp_grant),
      .PP_idle2_selected         (PP_idle2_selected),
      .PP_idle_selected          (PP_idle_selected),
      .PT_send_lreq              (PT_send_lreq),
      .PP_lreq_sent              (PP_lreq_sent),
      .PP_rx_data                (PP_rx_data),
      .PP_rx_charisk             (PP_rx_charisk),
      .PP_rx_valid               (PP_rx_valid),
      .PP_out_of_sync            (PP_out_of_sync),
      .PP_mode_1x                (PP_mode_1x),
      .PP_gttx_data              (PP_gttx_data),
      .PP_gttx_charisk           (PP_gttx_charisk),
      .PP_gttx_inhibit           (PP_gttx_inhibit),
      .GT_gtrx_data              (GT_gtrx_data),
      .GT_gtrx_charisk           (GT_gtrx_charisk),
      .GT_gtrx_chariscomma       (GT_gtrx_chariscomma),
      .GT_gtrx_disperr           (GT_gtrx_disperr),
      .GT_gtrx_notintable        (GT_gtrx_notintable),
      .PP_gtrx_chanbonden        (PP_gtrx_chanbonden),
      .GT_gtrx_chanisaligned     (GT_gtrx_chanisaligned),
      .GT_gtrx_reset_req         (GT_gtrx_reset_req),
      .PP_gtrx_reset             (PP_gtrx_reset),
      .GT_gtrx_reset_done        (GT_gtrx_reset_done),
      .PP_rx_lane_r              (PP_rx_lane_r),
      .PC_scram_disable          (PC_scram_disable),
      .PC_force_lane             (PC_force_lane),
      .PC_port_disable           (PC_port_disable),
      .PC_idle2_enable           (PC_idle2_enable),
      .PP_rx_scram_en            (PP_rx_scram_en),
      .PP_receiver_trained       (PP_receiver_trained),
      .PP_idle2_rcvd             (PP_idle2_rcvd),
      .PP_rx_lane_number         (PP_rx_lane_number),
      .PP_rx_port_width          (PP_rx_port_width),
      .PP_gt_decode_error        (PP_gt_decode_error),
      .PP_lane_sync              (PP_lane_sync),
//FIXCSF - CAL
// This is unsupported functionality, tie these to the appropriate ports
// once cs field command are allowed
      .PE_gttx_cmd               ({LINK_WIDTH{1'b0}}),
      .PE_gttx_tap_m1_cmd        ({LINK_WIDTH*2{1'b0}}),
      .PE_gttx_tap_p1_cmd        ({LINK_WIDTH*2{1'b0}}),
      .PE_gttx_reset_emphasis    ({LINK_WIDTH{1'b0}}),
      .PE_gttx_preset_emphasis   ({LINK_WIDTH{1'b0}}),
      .PE_gttx_tap_m1_status     ({LINK_WIDTH*2{1'b0}}),
      .PE_gttx_tap_p1_status     ({LINK_WIDTH*2{1'b0}}),
      .PE_gttx_ack               ({LINK_WIDTH{1'b0}}),
      .PE_gttx_nack              ({LINK_WIDTH{1'b0}}),
      .PP_gtrx_cmd               (),
      .PP_gtrx_tap_m1_cmd        (),
      .PP_gtrx_tap_p1_cmd        (),
      .PP_gtrx_reset_emphasis    (),
      .PP_gtrx_preset_emphasis   (),
      .PP_gtrx_tap_m1_status     (PP_gtrx_tap_m1_status),
      .PP_gtrx_tap_p1_status     (PP_gtrx_tap_p1_status),
      .PP_gtrx_ack               (),
      .PP_gtrx_nack              (),
      .PP_debug                  (PP_debug));
  // }}} End oplm_top inst

  // {{{ ollm_tx_top inst
  //--------------------------------------------
  srio_gen2_v4_1_16_ollm_tx_top
    #(.TCQ                       (TCQ),
      .LINK_WIDTH                (LINK_WIDTH),
      .GT_BYTES                  (GT_BYTES),
      .IDLE1                     (IDLE1),
      .IDLE2                     (IDLE2),
      .VC                        (VC),
      .SWITCH_MODE               (SWITCH_MODE),
      .SIM_TRAIN                 (SIM_TRAIN))
    ollm_tx_top_inst
     (.phy_clk                   (phy_clk),
      .phy_rst                   (phy_rst),
      .log_clk                   (log_clk),
      .log_rst                   (log_rst),
      .sim_train_en              (sim_train_en),
      .BT_phyt_tvalid            (BT_phyt_tvalid),
      .PT_phyt_tready            (PT_phyt_tready),
      .BT_phyt_tdata             (BT_phyt_tdata),
      .BT_phyt_tkeep             (BT_phyt_tkeep),
      .BT_phyt_tlast             (BT_phyt_tlast),
      .BT_phyt_tuser             (BT_phyt_tuser),
      .PT_phy_next_fm            (PT_phy_next_fm),
      .PT_sample_next_fm         (PT_sample_next_fm),
      .BT_tx_flow_control        (BT_tx_flow_control),
      .BR_phy_buf_stat           (BR_phy_buf_stat),
//FIXVC
//CAL - VCs not currently supported, need to link
//to the VC1 status when integrated, for now
//it can be the VC0 buf_stat
      .BR_phy_buf_stat_vc1       (BR_phy_buf_stat),
      .PP_port_initialized       (PP_port_initialized),
      .PP_mode_1x                (PP_mode_1x),
      .PP_idle2_selected         (PP_idle2_selected),
      .PT_tx_data                (PT_tx_data),
      .PT_tx_charisk             (PT_tx_charisk),
      .PT_tx_valid               (PT_tx_valid),
      .PT_tx_early_valid         (PT_tx_early_valid),
      .PT_tx_early_lreq          (PT_tx_early_lreq),
      .PP_ccomp_req              (PP_ccomp_req),
      .PT_ccomp_grant            (PT_ccomp_grant),
      .PT_send_lreq              (PT_send_lreq),
      .PP_lreq_sent              (PP_lreq_sent),
      .PC_send_lreq              (PC_send_lreq),
      .PC_lreq_cmd               (PC_lreq_cmd),
      .PC_load_ackids            (PC_load_ackids),
      .PC_load_nextpkt           (PC_load_nextpkt),
      .PC_next_fm                (PC_next_fm),
      .PC_vc_en                  (PC_vc_en),
//FIXVC
//CAL - VCs not currently supported, need to link to the
//PC when integrated.
      .PC_vc1_refresh_int        (8'h00),
      .PR_link_initialized       (PR_link_initialized),
      .PT_sent_init_cs           (PT_sent_init_cs),
      .PR_rewind                 (PR_rewind),
      .PT_phy_rewind             (PT_phy_rewind),
      .PR_phy_last_ack           (PR_phy_last_ack),
      .PR_send_rfr               (PR_send_rfr),
      .PT_rfr_sent               (PT_rfr_sent),
      .PR_send_lreq              (PR_send_lreq),
      .PT_lreq_sent              (PT_lreq_sent),
      .PR_send_pna               (PR_send_pna),
      .PT_pna_sent               (PT_pna_sent),
      .PR_send_pr                (PR_send_pr),
      .PT_pr_sent                (PT_pr_sent),
      .PR_send_lresp             (PR_send_lresp),
      .PT_lresp_sent             (PT_lresp_sent),
      .PR_last_good_pkt          (PR_last_good_pkt),
      .PR_cause                  (PR_cause),
      .PR_port_stat              (PR_port_stat),
      .PT_switch_crc_err         (PT_switch_crc_err),
      .PR_output_error_stop      (PR_output_error_stop),
      .PR_rcvd_error_free_status (PR_rcvd_error_free_status),
      .UG_phy_mce                (UG_phy_mce),
      .UG_phy_link_reset         (UG_phy_link_reset),
      .PT_debug                  (PT_debug));
  // }}} end ollm_tx_top inst

  // {{{ ollm_rx_top instantiation
  //--------------------------------------------
  srio_gen2_v4_1_16_ollm_rx_top
    #(.TCQ                       (TCQ),
      .IDLE1                     (IDLE1),
      .IDLE2                     (IDLE2),
      .MODE_XG                   (MODE_XG),
      .VC                        (VC),
      .SWITCH_MODE               (SWITCH_MODE),
      .RETRY                     (RETRY),
      .TARGET_DS                 (TARGET_DS),
      .LINK_REQUESTS             (LINK_REQUESTS),
      .VC1_CT                    (VC1_CT),
      .LINK_WIDTH                (LINK_WIDTH))

    ollm_rx_top_inst
     (.phy_clk                   (phy_clk),
      .phy_rst                   (phy_rst),
      .log_clk                   (log_clk),
      .log_rst                   (log_rst),
      .gt_pcs_clk                (gt_pcs_clk),
      .PR_phy_rcvd_mce           (PR_phy_rcvd_mce),
      .PR_phy_rcvd_link_reset    (PR_phy_rcvd_link_reset),
      .PR_debug                  (PR_debug),

      .PP_rx_data                (PP_rx_data),
      .PP_rx_charisk             (PP_rx_charisk),
      .PP_rx_valid               (PP_rx_valid),
      .PP_idle2_selected         (PP_idle2_selected),
      .PP_out_of_sync            (PP_out_of_sync),
      .PP_port_initialized       (PP_port_initialized),
      .PP_mode_1x                (PP_mode_1x),
      .PP_gt_decode_error        (PP_gt_decode_error),

      .PR_phyr_tvalid            (PR_phyr_tvalid),
      .BR_phyr_tready            (BR_phyr_tready),
      .PR_phyr_tdata             (PR_phyr_tdata),
      .PR_phyr_tkeep             (PR_phyr_tkeep),
      .PR_phyr_tlast             (PR_phyr_tlast),
      .PR_phyr_tuser             (PR_phyr_tuser),
      .BR_phy_buf_stat           (BR_phy_buf_stat),

      .PT_sent_init_cs           (PT_sent_init_cs),
      .PR_link_initialized       (PR_link_initialized),
      .PR_rewind                 (PR_rewind),
      .PR_phy_last_ack           (PR_phy_last_ack),
      .PT_phy_next_fm            (PT_phy_next_fm),
      .PR_phy_rcvd_buf_stat      (PR_phy_rcvd_buf_stat),
      .PR_send_rfr               (PR_send_rfr),
      .PT_rfr_sent               (PT_rfr_sent),
      .PR_send_lreq              (PR_send_lreq),
      .PT_lreq_sent              (PT_lreq_sent),
      .PR_send_pna               (PR_send_pna),
      .PT_pna_sent               (PT_pna_sent),
      .PR_send_pr                (PR_send_pr),
      .PT_pr_sent                (PT_pr_sent),
      .PR_send_lresp             (PR_send_lresp),
      .PT_lresp_sent             (PT_lresp_sent),
      .PR_cause                  (PR_cause),
      .PR_port_stat              (PR_port_stat),
      .PR_last_good_pkt          (PR_last_good_pkt),
      .PR_output_retry_stop      (PR_output_retry_stop),
      .PR_output_error_stop      (PR_output_error_stop),
      .PR_port_error             (PR_port_error),
      .PR_input_retry_stop       (PR_input_retry_stop),
      .PR_input_error_stop       (PR_input_error_stop),
      .PR_rcvd_error_free_status (PR_rcvd_error_free_status),
      .PT_sample_next_fm         (PT_sample_next_fm),

      .PR_next_rcvd_pkt          (PR_next_rcvd_pkt),
      .PC_last_ack               (PC_last_ack),
      .PC_load_ackids            (PC_load_ackids),
      .PC_load_nextpkt           (PC_load_nextpkt),
      .PC_send_lreq              (PC_send_lreq),
      .PC_lreq_cmd               (PC_lreq_cmd),
      .PC_link_timeout           (PC_link_timeout),
      .PC_clr_port_error         (PC_clr_port_error),
      .PC_input_maint_only       (PC_input_maint_only),
      .PC_error_disable          (PC_error_disable),
      .PC_vc_ct                  (PC_vc_ct),
      .PC_vc_en                  (PC_vc_en),
      .PR_rcvd_lresp             (PR_rcvd_lresp),
      .PR_ackid_status           (PR_ackid_status),
      .PR_rcvd_port_stat         (PR_rcvd_port_stat),
      .PC_next_rcvd_pkt          (PC_next_rcvd_pkt),
      .PR_rcvd_pa_or_pna         (PR_rcvd_pa_or_pna));
  // }}} End ollm_rx_top inst

  // {{{ phy_cfg_top instantiation
  //--------------------------------------------
  srio_gen2_v4_1_16_phy_cfg_top
    #(.TCQ                       (TCQ),
      .PHY_EF_PTR                (PHY_EF_PTR),
      .LANE_EF_PTR               (LANE_EF_PTR),
      .VC_EF_PTR                 (VC_EF_PTR),
      .USER_EF_PTR               (USER_EF_PTR),
      .LINK_TIMEOUT              (LINK_TIMEOUT),
      .PORT_TIMEOUT              (PORT_TIMEOUT),
      .SW_CSR                    (SW_CSR),
      .VC                        (VC),
      .VC1_CT                    (VC1_CT),
      .IS_HOST                   (IS_HOST),
      .MASTER_EN                 (MASTER_EN),
      .DISCOVERED                (DISCOVERED),
      .IDLE1                     (IDLE1),
      .IDLE2                     (IDLE2),
      .MODE_XG                   (MODE_XG),
      .GT_BYTES                  (GT_BYTES),
      .LINK_WIDTH                (LINK_WIDTH))
    phy_cfg_top_inst
     (.phy_clk                   (phy_clk),
      .phy_rst                   (phy_rst),
      .gt_pcs_clk                (gt_pcs_clk),
      .gt_pcs_rst                (gt_pcs_rst),
      .cfg_clk                   (cfg_clk),
      .cfg_rst                   (cfg_rst),
      .PC_port_timeout           (PC_port_timeout),
      .PC_srio_host              (PC_srio_host),
      .PC_maint_only             (PC_maint_only),
      .PC_master_enable          (PC_master_enable),
      .BT_tx_flow_control        (BT_tx_flow_control),
      .PT_phy_next_fm            (PT_phy_next_fm),
      .PC_next_fm                (PC_next_fm),
      .PC_lreq_cmd               (PC_lreq_cmd),
      .PC_send_lreq              (PC_send_lreq),
      .PC_load_ackids            (PC_load_ackids),
      .PC_load_nextpkt           (PC_load_nextpkt),
      .PR_phy_last_ack           (PR_phy_last_ack),
      .PR_next_rcvd_pkt          (PR_next_rcvd_pkt),
      .PR_rcvd_lresp             (PR_rcvd_lresp),
      .PR_ackid_status           (PR_ackid_status),
      .PR_rcvd_port_stat         (PR_rcvd_port_stat),
      .PR_output_retry_stop      (PR_output_retry_stop),
      .PR_output_error_stop      (PR_output_error_stop),
      .PR_input_retry_stop       (PR_input_retry_stop),
      .PR_input_error_stop       (PR_input_error_stop),
      .PR_rcvd_pa_or_pna         (PR_rcvd_pa_or_pna),
      .PR_port_error             (PR_port_error),
      .PC_next_rcvd_pkt          (PC_next_rcvd_pkt),
      .PC_last_ack               (PC_last_ack),
      .PC_link_timeout           (PC_link_timeout),
      .PC_vc_ct                  (PC_vc_ct),
      .PC_vc_en                  (PC_vc_en),
      .PC_input_maint_only       (PC_input_maint_only),
      .PC_error_disable          (PC_error_disable),
      .PC_clr_port_error         (PC_clr_port_error),
      .PP_idle_selected          (PP_idle_selected),
      .PP_idle2_selected         (PP_idle2_selected),
      .PP_mode_1x                (PP_mode_1x),
      .PP_port_initialized       (PP_port_initialized),
      .PP_rx_lane_r              (PP_rx_lane_r),
      .PP_gtrx_tap_m1_status     (PP_gtrx_tap_m1_status),
      .PP_gtrx_tap_p1_status     (PP_gtrx_tap_p1_status),
      .PP_rx_scram_en            (PP_rx_scram_en),
      .PP_receiver_trained       (PP_receiver_trained),
      .PP_idle2_rcvd             (PP_idle2_rcvd),
      .PP_rx_lane_number         (PP_rx_lane_number),
      .PP_rx_port_width          (PP_rx_port_width),
      .PP_gt_decode_error        (PP_gt_decode_error),
      .PP_lane_sync              (PP_lane_sync),
      .PC_force_lane             (PC_force_lane),
      .PC_scram_disable          (PC_scram_disable),
      .PC_port_disable           (PC_port_disable),
      .PC_idle2_enable           (PC_idle2_enable),
      .CF_cfgp_awvalid           (CF_cfgp_awvalid),
      .PC_cfgp_awready           (PC_cfgp_awready),
      .CF_cfgp_awaddr            (CF_cfgp_awaddr),
      .CF_cfgp_wvalid            (CF_cfgp_wvalid),
      .PC_cfgp_wready            (PC_cfgp_wready),
      .CF_cfgp_wdata             (CF_cfgp_wdata),
      .CF_cfgp_wstrb             (CF_cfgp_wstrb),
      .PC_cfgp_bvalid            (PC_cfgp_bvalid),
      .CF_cfgp_bready            (CF_cfgp_bready),
      .CF_cfgp_arvalid           (CF_cfgp_arvalid),
      .PC_cfgp_arready           (PC_cfgp_arready),
      .CF_cfgp_araddr            (CF_cfgp_araddr),
      .PC_cfgp_rvalid            (PC_cfgp_rvalid),
      .CF_cfgp_rready            (CF_cfgp_rready),
      .PC_cfgp_rdata             (PC_cfgp_rdata));
  // }}} End phy_cfg_top inst

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/phy/ollm_tx/srio_gen2_v4_1_16_ollm_tx_top.v#1 $
//----------------------------------------------------------------------
//
// OLLM_TX_TOP
// Description:
// This module instantiates all the submodules of the OLLM TX design
//
// Hierarchy:
// PHY_TOP
//    |___OLLM_TX_TOP <-- this module
//             |_____OLLM_TX_READY_GEN
//             |_____OLLM_TX_BUF
//             |_____OLLM_TX_PKT_ASSEMBLY
//             |_____OLLM_TX_CS_GEN
//             |_____OLLM_TX_DATA_MUX
//             |_____OLLM_TX_OPLM
// ---------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_ollm_tx_top
  #(
    parameter TCQ         = 100,
    parameter LINK_WIDTH  = 1,    // Generated Link Width {1, 2, 4}
    parameter GT_BYTES    = 4,    // Bytes per cycle on the GT Interface
    parameter IDLE1       = 1,    // Include the IDLE1 Sequence {0,1}
    parameter IDLE2       = 0,    // Include the IDLE2 Sequence {0,1}
    parameter VC          = 0,    // Highest numbered VC supported {0,1}
    parameter SWITCH_MODE = 0,    // If the core support Switch Mode
    parameter SIM_TRAIN   = 0)    // {0: FULL, 1: DIVIDED, 3: TRAINED}
  (
    // {{{ Port Declarations
    // System Signals
    input             phy_clk,                  // PHY interface clock
    input             phy_rst,                  // Reset for PHY clock Domain
    input             log_clk,                  // LOG interface clock
    input             log_rst,                  // Reset for LOG clock Domain
    input             sim_train_en,             // Enable the SIM_TRAIN parameter

    //TX Buffer Interface Signals
    input             BT_phyt_tvalid,           // Valid data indicator
    output            PT_phyt_tready,           // Destination Ready
    input  [63:0]     BT_phyt_tdata,            // Packet for transfer
    input  [7:0]      BT_phyt_tkeep,            // Byte Enable for transferred packet
    input             BT_phyt_tlast,            // Last DW of incoming packet
    input  [7:0]      BT_phyt_tuser,            // {1'b0, SKIP_CRC, 2'h00, VC[1:0], CRF, SRC_DSC}
    output [5:0]      PT_phy_next_fm,           // Next packets AckID
    output            PT_sample_next_fm,        // Indicates to the ollm rx to sample the next fm
                                                //  value in a rewind scenario.
    output            PT_phy_rewind,            // Holds PR_rewind high as long as we
                                                //  are killing a packet
    input             BT_tx_flow_control,       // Flow Control Mode of the TX Buffer

    //RX Buffer Interface Signals
    input  [5:0]      BR_phy_buf_stat,          // VC0 status from the RX buffer
    input  [5:0]      BR_phy_buf_stat_vc1,      // VC1 status from the RX buffer

    //OPLM TX Interface Signals
    input             PP_port_initialized,      // Indicates port is initialized
    input             PP_mode_1x,               // Indicates the link trained down to 1x
    input             PP_idle2_selected,        // Indicated the operating idle mode
    output [63:0]     PT_tx_data,               // Transmit data
    output [7:0]      PT_tx_charisk,            // Indicates which bytes  are K characters
    output [1:0]      PT_tx_valid,              // Indicates valid words
    output [1:0]      PT_tx_early_valid,        // Indicates valid words upcoming in two cycles
    output            PT_tx_early_lreq,         // Indicates an lreq upcoming in two cycles
    input             PP_ccomp_req,             // Request break for clock compensation sequence
    output            PT_ccomp_grant,           // Insert clock compensation at next invalid
    output            PT_send_lreq,             // Indicates the data on PT_tx_data is a LREQ
    input             PP_lreq_sent,             // Indicates the LREQ SYNC SEQ was sent

    //PHY Config Interface Signals
    input             PC_send_lreq,             // Send a Link Request Input Status CS
    input  [2:0]      PC_lreq_cmd,              // Command information for PC_send_lreq
    input             PC_load_ackids,           // Indication to load PC_next_fm into phy_next_fm
    input             PC_load_nextpkt,          // Indicated when a new ackid is loaded in the ollm rx
    input  [5:0]      PC_next_fm,               // Value to load into phy_next_fm when
                                                //  PC_load_ackids is asserted
    input             PC_vc_en,                 // Enable VC1
    input  [7:0]      PC_vc1_refresh_int,       // The Refresh Interval for VC1

    //OLLM RX Interface Signals
    input             PR_link_initialized,      // Indicates the link is initialized
    output            PT_sent_init_cs,          // Indicates the link init seq. was sent

    input             PR_rewind,                // Indicates error or retry condition and the
                                                //  next_fm must be updated
    input  [5:0]      PR_phy_last_ack,          // Last PA received by the PHY core

    input             PR_send_rfr,              // Send an RFR control symbol (Request)
    output            PT_rfr_sent,              // Sent RFR (Grant)
    input             PR_send_lreq,             // Send a Link Request Input Status
    output            PT_lreq_sent,             // Sent Link Request Input Status
    input             PR_send_pna,              // Send a PNA control symbol
    output            PT_pna_sent,              // Sent PNA
    input             PR_send_pr,               // Send a PR control symbol
    output            PT_pr_sent,               // Sent PR
    input             PR_send_lresp,            // Send a Link Response Control Symbol
    output            PT_lresp_sent,            // Sent Link Response

    input  [5:0]      PR_last_good_pkt,         // Last PA to send
    input  [4:0]      PR_cause,                 // Last cause for a PNA to send
    input  [4:0]      PR_port_stat,             // Current port status
    output            PT_switch_crc_err,        // A crc error was detected in switch mode
    input             PR_output_error_stop,     // The OLLM RX is in the output error stopped state
    input             PR_rcvd_error_free_status,// Indicates when an error free status cs
                                                //  is recieved from the link partner
    //User Interface Signals
    input             UG_phy_mce,               // Send MCE control symbol
    input             UG_phy_link_reset,        // Send link reset control symbols

    //Debug Interface
    output [63:0]     PT_debug                  // OLLM TX debug bus, should include useful
                                                //  signals for HW debug
    // }}} end Port Declarations
  );

  // {{{ Wire Declarations
  // Throughout this code the three letter prefixs indicate the following:
  // PTB = OLLM TX Buffer
  // PTA = OLLM TX Assembly
  // PTS = OLLM TX Symbols
  // PTM = OLLM TX Mux
  // PTP = OLLM TX OPLM
  // PTR = OLLM TX Ready Gen

  //Signals from packet stack to tx buf if
  wire          BT_phyt_tvalid_stack;
  wire          PT_phyt_tready_stack;
  wire [63:0]   BT_phyt_tdata_stack;
  wire [7:0]    BT_phyt_tkeep_stack;
  wire          BT_phyt_tlast_stack;
  wire [7:0]    BT_phyt_tuser_stack;
  wire          PT_phy_rewind_int;

  //Signals from tx buf if to packet assembly
  wire  [5:0]   PTB_next_fm;
  wire          PTB_sop;
  wire          PTB_eop;
  wire          PTB_src_disc; // CR 800810, stomp
  wire          PTB_valid;
  wire          PTB_valid_d;
  wire  [63:0]  PTB_data;
  wire  [3:0]   PTB_keep;
  wire          PTB_vc;
  wire          PTB_crf;
  wire          PTB_in_packet;
  wire          PTB_skip_final_crc;
  wire  [15:0]  PTB_crc64;
  wire  [15:0]  PTB_crc48;
  wire  [15:0]  PTB_crc32;
  wire  [15:0]  PTB_crc16;
  wire          PTB_insert_mid_crc;
  wire          PTB_mid_crc_inserted;

  // Signals from the tx buf if to the cs generator
  wire          PTB_sop_d;
  wire          PTB_link_reset;

  //Signals from packet assembly to the data mux
  wire          PTA_sop;
  wire          PTA_eop;
  wire          PTA_in_packet;
  wire          PTA_in_packet_d;
  wire [63:0]   PTA_data;
  wire [1:0]    PTA_valid;
  wire [1:0]    PTA_valid_d;
  wire          PTA_eop_d;

  //Signals from the cs gen block to the data mux
  wire [63:0]   PTS_data;
  wire [1:0]    PTS_valid;
  wire          PTS_lreq;
  wire          PTS_embed_cs;
  wire [7:0]    PTS_charisk;
  wire          PTS_sop;
  wire          PTS_eop;
  wire          PTS_stall;

  //Signals from the data mux to the oplm interface
  wire [63:0]   PTM_data;
  wire [1:0]    PTM_valid;
  wire [7:0]    PTM_charisk;
  wire          PTM_send_lreq;

  //Signals from the Ready generator to the other modules
  wire          PTR_ptp_advance;
  wire          PTR_ptm_advance;
  wire          PTR_pta_advance;
  wire          PTR_pts_advance;
  wire          PTR_ptb_advance;

  //Stall Signals to the ready generator
  wire          PTB_stall;
  wire          PTP_stall;
  wire          PTM_pta_stall;
  wire          PTM_pts_stall;
  wire          PTA_stall;

  // Signals to the debug bus
  wire          PTS_mce_sent;
  wire          PTS_pa_sent;

  // Set the debug bus
  assign PT_debug[0] = PT_rfr_sent;
  assign PT_debug[1] = PT_lreq_sent;
  assign PT_debug[2] = PT_pna_sent;
  assign PT_debug[3] = PT_pr_sent;
  assign PT_debug[4] = PT_lresp_sent;
  assign PT_debug[5] = PTS_mce_sent;
  assign PT_debug[6] = PTS_pa_sent;       // A PA is sent for each cycle this is asserted
  assign PT_debug[7] = PT_sent_init_cs;   // Asserted when all 15-Status CSs have been sent for link init
  assign PT_debug[8] = PC_send_lreq;      // Asserted until a LREQ is sent
  assign PT_debug[9] = PTB_link_reset;    // Asserted as long as LREQ/resets must stream,
                                          // may have delayed assertion until its safe for
                                          // the core to stream these
  assign PT_debug[63:10] = 54'b0;
  // }}} end Wire Declarations


  // {{{ ollm_tx_pkt_stack inst
  //--------------------------------------------
  srio_gen2_v4_1_16_ollm_tx_pkt_stack
    #(.TCQ                       (TCQ),
      .BYPASS                    (0))
    ollm_tx_pkt_stack_inst
     (.phy_clk                   (phy_clk),
      .phy_rst                   (phy_rst),

      .BT_phyt_tvalid            (BT_phyt_tvalid),
      .PT_phyt_tready            (PT_phyt_tready),
      .BT_phyt_tdata             (BT_phyt_tdata),
      .BT_phyt_tkeep             (BT_phyt_tkeep),
      .BT_phyt_tlast             (BT_phyt_tlast),
      .BT_phyt_tuser             (BT_phyt_tuser),

      .BT_phyt_tvalid_stack      (BT_phyt_tvalid_stack),
      .PT_phyt_tready_stack      (PT_phyt_tready_stack),
      .BT_phyt_tdata_stack       (BT_phyt_tdata_stack),
      .BT_phyt_tkeep_stack       (BT_phyt_tkeep_stack),
      .BT_phyt_tlast_stack       (BT_phyt_tlast_stack),
      .BT_phyt_tuser_stack       (BT_phyt_tuser_stack),

      .PT_phy_rewind             (PT_phy_rewind),
      .PT_phy_rewind_int         (PT_phy_rewind_int));

  // }}} end ollm_tx_pkt_stack inst

  // {{{ ollm_tx_buf inst
  //--------------------------------------------
  srio_gen2_v4_1_16_ollm_tx_buf
    #(.TCQ                       (TCQ),
      .IDLE1                     (IDLE1),
      .IDLE2                     (IDLE2),
      .SWITCH_MODE               (SWITCH_MODE))
    ollm_tx_buf_inst
     (.phy_clk                   (phy_clk),
      .phy_rst                   (phy_rst),
      .BT_phyt_tvalid            (BT_phyt_tvalid_stack),
      .PT_phyt_tready            (PT_phyt_tready_stack),
      .BT_phyt_tdata             (BT_phyt_tdata_stack),
      .BT_phyt_tkeep             (BT_phyt_tkeep_stack),
      .BT_phyt_tlast             (BT_phyt_tlast_stack),
      .BT_phyt_tuser             (BT_phyt_tuser_stack),
      .PTB_phy_next_fm           (PT_phy_next_fm),
      .PTB_sample_next_fm        (PT_sample_next_fm),
      .UG_phy_link_reset         (UG_phy_link_reset),
      .PTB_next_fm               (PTB_next_fm),
      .PTB_sop_d                 (PTB_sop_d),
      .PTB_sop                   (PTB_sop),
      .PTB_eop                   (PTB_eop),
      .PTB_src_disc              (PTB_src_disc), // cr 800810, stomp
      .PTB_valid                 (PTB_valid),
      .PTB_valid_d               (PTB_valid_d),
      .PTB_in_packet             (PTB_in_packet),
      .PTB_data                  (PTB_data),
      .PTB_keep                  (PTB_keep),
      .PTB_vc                    (PTB_vc),
      .PTB_crf                   (PTB_crf),
      .PTB_skip_final_crc        (PTB_skip_final_crc),
      .PTB_crc64                 (PTB_crc64),
      .PTB_crc48                 (PTB_crc48),
      .PTB_crc32                 (PTB_crc32),
      .PTB_crc16                 (PTB_crc16),
      .PTB_insert_mid_crc        (PTB_insert_mid_crc),
      .PTB_mid_crc_inserted      (PTB_mid_crc_inserted),
      .PTS_lreq_sent             (PT_lreq_sent),
      .PTS_rfr_sent              (PT_rfr_sent),
      .PR_send_rfr               (PR_send_rfr),
      .PR_send_lreq              (PR_send_lreq),
      .PTB_link_reset            (PTB_link_reset),
      .PR_rewind                 (PR_rewind),
      .PR_link_initialized       (PR_link_initialized),
      .PTB_phy_rewind            (PT_phy_rewind_int),
      .PR_phy_last_ack           (PR_phy_last_ack),
      .PP_port_initialized       (PP_port_initialized),
      .PP_idle2_selected         (PP_idle2_selected),
      .PC_load_ackids            (PC_load_ackids),
      .PC_next_fm                (PC_next_fm),
      .PTB_stall                 (PTB_stall),
      .PTR_ptb_advance           (PTR_ptb_advance));

  // }}} end ollm_tx_buf inst

  // {{{ ollm_tx_pkt_assembly inst
  //--------------------------------------------
  srio_gen2_v4_1_16_ollm_tx_pkt_assembly
    #(.TCQ                       (TCQ),
      .IDLE2                     (IDLE2),
      .SWITCH_MODE               (SWITCH_MODE))
    ollm_tx_pkt_assembly_inst
     (.phy_clk                   (phy_clk),
      .phy_rst                   (phy_rst),
      .PT_switch_crc_err         (PT_switch_crc_err),
      .PTB_sop                   (PTB_sop),
      .PTB_eop                   (PTB_eop),
      .PTB_valid                 (PTB_valid),
      .PTB_valid_d               (PTB_valid_d),
      .PTB_data                  (PTB_data),
      .PTB_keep                  (PTB_keep),
      .PTB_vc                    (PTB_vc),
      .PTB_crf                   (PTB_crf),
      .PTB_skip_final_crc        (PTB_skip_final_crc),
      .PTB_in_packet             (PTB_in_packet),
      .PTB_crc64                 (PTB_crc64),
      .PTB_crc48                 (PTB_crc48),
      .PTB_crc32                 (PTB_crc32),
      .PTB_crc16                 (PTB_crc16),
      .PTB_insert_mid_crc        (PTB_insert_mid_crc),
      .PTB_mid_crc_inserted      (PTB_mid_crc_inserted),
      .PTB_next_fm               (PTB_next_fm),
      .PTA_data                  (PTA_data),
      .PTA_valid_d               (PTA_valid_d),
      .PTA_valid                 (PTA_valid),
      .PTA_sop                   (PTA_sop),
      .PTA_eop_d                 (PTA_eop_d),
      .PTA_eop                   (PTA_eop),
      .PTA_in_packet             (PTA_in_packet),
      .PTA_in_packet_d           (PTA_in_packet_d),
      .PP_idle2_selected         (PP_idle2_selected),
      .PTA_stall                 (PTA_stall),
      .PTR_pta_advance           (PTR_pta_advance));
  // }}} end ollm_tx_pkt_assembly inst

  // {{{ ollm_tx_cs_gen inst
  //--------------------------------------------
  srio_gen2_v4_1_16_ollm_tx_cs_gen
    #(.TCQ                       (TCQ),
      .LINK_WIDTH                (LINK_WIDTH),
      .GT_BYTES                  (GT_BYTES),
      .IDLE1                     (IDLE1),
      .IDLE2                     (IDLE2),
      .VC                        (VC),
      .SIM_TRAIN                 (SIM_TRAIN))
    ollm_tx_cs_gen_inst
     (.phy_clk                   (phy_clk),
      .phy_rst                   (phy_rst),
      .log_clk                   (log_clk),
      .log_rst                   (log_rst),
      .sim_train_en              (sim_train_en),
      .BT_tx_flow_control        (BT_tx_flow_control),
      .BR_phy_buf_stat           (BR_phy_buf_stat),
      .BR_phy_buf_stat_vc1       (BR_phy_buf_stat_vc1),
      .PP_port_initialized       (PP_port_initialized),
      .PP_mode_1x                (PP_mode_1x),
      .PP_idle2_selected         (PP_idle2_selected),
      .PP_ccomp_req              (PP_ccomp_req),
      .PT_ccomp_grant            (PT_ccomp_grant),
      .PC_send_lreq              (PC_send_lreq),
      .PC_lreq_cmd               (PC_lreq_cmd),
      .PC_vc_en                  (PC_vc_en),
      .PC_vc1_refresh_int        (PC_vc1_refresh_int),
      .PC_load_nextpkt           (PC_load_nextpkt),
      .PTS_sent_init_cs          (PT_sent_init_cs),
      .PR_send_rfr               (PR_send_rfr),
      .PTS_rfr_sent              (PT_rfr_sent),
      .PR_send_lreq              (PR_send_lreq),
      .PTS_lreq_sent             (PT_lreq_sent),
      .PR_send_pna               (PR_send_pna),
      .PTS_pna_sent              (PT_pna_sent),
      .PR_send_pr                (PR_send_pr),
      .PTS_pr_sent               (PT_pr_sent),
      .PR_send_lresp             (PR_send_lresp),
      .PTS_lresp_sent            (PT_lresp_sent),
      .PR_last_good_pkt          (PR_last_good_pkt),
      .PR_cause                  (PR_cause),
      .PR_port_stat              (PR_port_stat),
      .PR_link_initialized       (PR_link_initialized),
      .PR_output_error_stop      (PR_output_error_stop),
      .PR_rcvd_error_free_status (PR_rcvd_error_free_status),
      .UG_phy_mce                (UG_phy_mce),
      .PTB_sop_d                 (PTB_sop_d),
      .PTB_sop                   (PTB_sop),
      .PTB_src_disc              (PTB_src_disc), // cr 800810, stomp
      .PTB_eop                   (PTB_eop),
      .PTB_next_fm               (PTB_next_fm),
      .PTR_ptb_advance           (PTR_ptb_advance),
      .PTB_in_packet             (PTB_in_packet),
      .PTB_link_reset            (PTB_link_reset),
      .PTA_in_packet             (PTA_in_packet),
      .PTA_valid_d               (PTA_valid_d),
      .PTA_eop                   (PTA_eop),
      .PTR_pta_advance           (PTR_pta_advance),
      .PTS_data                  (PTS_data),
      .PTS_valid                 (PTS_valid),
      .PTS_lreq                  (PTS_lreq),
      .PTS_embed_cs              (PTS_embed_cs),
      .PTS_charisk               (PTS_charisk),
      .PTS_sop                   (PTS_sop),
      .PTS_eop                   (PTS_eop),
      .PTS_stall                 (PTS_stall),
      .PTR_pts_advance           (PTR_pts_advance),
      .PTS_mce_sent              (PTS_mce_sent),
      .PTS_pa_sent               (PTS_pa_sent));
  // }}} end ollm_tx_cs_gen inst

  // {{{ ollm_tx_data_mux inst
  //--------------------------------------------
  srio_gen2_v4_1_16_ollm_tx_data_mux
    #(.TCQ                       (TCQ))
    ollm_tx_data_mux_inst
     (.phy_clk                   (phy_clk),
      .phy_rst                   (phy_rst),
      .PT_phy_rewind             (PT_phy_rewind_int),
      .PTA_data                  (PTA_data),
      .PTA_valid_d               (PTA_valid_d),
      .PTA_valid                 (PTA_valid),
      .PTA_sop                   (PTA_sop),
      .PTA_eop_d                 (PTA_eop_d),
      .PTA_eop                   (PTA_eop),
      .PTA_in_packet             (PTA_in_packet),
      .PTA_in_packet_d           (PTA_in_packet_d),
      .PTS_data                  (PTS_data),
      .PTS_valid                 (PTS_valid),
      .PTS_lreq                  (PTS_lreq),
      .PTS_embed_cs              (PTS_embed_cs),
      .PTS_charisk               (PTS_charisk),
      .PTS_sop                   (PTS_sop),
      .PTS_eop                   (PTS_eop),
      .PR_link_initialized       (PR_link_initialized),
      .PP_ccomp_req              (PP_ccomp_req),
      .PP_idle2_selected         (PP_idle2_selected),
      .PTM_data                  (PTM_data),
      .PTM_valid                 (PTM_valid),
      .PTM_charisk               (PTM_charisk),
      .PTM_send_lreq             (PTM_send_lreq),
      .PTM_tx_early_valid        (PT_tx_early_valid),
      .PTM_tx_early_lreq         (PT_tx_early_lreq),
      .PTM_pta_stall             (PTM_pta_stall),
      .PTM_pts_stall             (PTM_pts_stall),
      .PTR_pta_advance           (PTR_pta_advance),
      .PTR_pts_advance           (PTR_pts_advance),
      .PTR_ptm_advance           (PTR_ptm_advance));

  // }}} end ollm_tx_data_mux inst

  // {{{ ollm_tx_oplm inst
  //--------------------------------------------
  srio_gen2_v4_1_16_ollm_tx_oplm
    #(.TCQ                       (TCQ))
    ollm_tx_oplm_inst
     (.phy_clk                   (phy_clk),
      .phy_rst                   (phy_rst),
      .PTM_data                  (PTM_data),
      .PTM_valid                 (PTM_valid),
      .PTM_charisk               (PTM_charisk),
      .PTM_send_lreq             (PTM_send_lreq),
      .PTP_tx_data               (PT_tx_data),
      .PTP_tx_charisk            (PT_tx_charisk),
      .PTP_tx_valid              (PT_tx_valid),
      .PP_ccomp_req              (PP_ccomp_req),
      .PTP_ccomp_grant           (PT_ccomp_grant),
      .PTP_send_lreq             (PT_send_lreq),
      .PP_lreq_sent              (PP_lreq_sent),
      .PTP_stall                 (PTP_stall),
      .PTR_ptp_advance           (PTR_ptp_advance));
  // }}} end ollm_tx_top inst

  // {{{ ollm_tx_ready_gen inst
  //--------------------------------------------
  srio_gen2_v4_1_16_ollm_tx_ready_gen
    #(.TCQ    (TCQ))
    ollm_tx_ready_gen_inst
      (.phy_clk             (phy_clk),
       .phy_rst             (phy_rst),
       .PTR_phyt_tready     (PT_phyt_tready_stack),
       .PTB_stall           (PTB_stall),
       .PTR_ptb_advance     (PTR_ptb_advance),
       .PTP_stall           (PTP_stall),
       .PTR_ptp_advance     (PTR_ptp_advance),
       .PTM_pta_stall       (PTM_pta_stall),
       .PTM_pts_stall       (PTM_pts_stall),
       .PTR_ptm_advance     (PTR_ptm_advance),
       .PTA_in_packet       (PTA_in_packet),
       .PTA_stall           (PTA_stall),
       .PTR_pta_advance     (PTR_pta_advance),
       .PTS_stall           (PTS_stall),
       .PTR_pts_advance     (PTR_pts_advance));
   // }}} end ollm_tx_ready_gen inst


endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/phy/ollm_tx/srio_gen2_v4_1_16_ollm_tx_top.v#3 $
//----------------------------------------------------------------------
//
// OLLM_TX_TOP
// Description:
// This module plugs in between the buffer tx and the OLLM TX
// This was created afterwards to improve some noted performance problems and
// can be removed to save resources at the expence of performance
//
// Hierarchy:
// PHY_TOP
//    |___OLLM_TX_TOP <-- this module
//             |_____OLLM_TX_READY_GEN
//             |_____OLLM_TX_PKT_STACK
//             |_____OLLM_TX_BUF
//             |_____OLLM_TX_PKT_ASSEMBLY
//             |_____OLLM_TX_CS_GEN
//             |_____OLLM_TX_DATA_MUX
//             |_____OLLM_TX_OPLM
// ---------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_ollm_tx_pkt_stack
  #(
    parameter TCQ         = 100,
    parameter BYPASS      = 0)  // When set, directly wire ins to outs
  (
    // {{{ Port Declarations
    // System Signals
    input             phy_clk,                  // PHY interface clock
    input             phy_rst,                  // Reset for PHY clock Domain

    // TX Buffer Interface Signals
    input             BT_phyt_tvalid,           // Valid data indicator
    output            PT_phyt_tready,           // Destination Ready
    input  [63:0]     BT_phyt_tdata,            // Packet for transfer
    input  [7:0]      BT_phyt_tkeep,            // Byte Enable for transferred packet
    input             BT_phyt_tlast,            // Last DW of incoming packet
    input  [7:0]      BT_phyt_tuser,            // {1'b0, SKIP_CRC, 2'h00, VC[1:0], CRF, SRC_DSC} 


    // OLLM TX internal signals
    output            BT_phyt_tvalid_stack,     // Valid data indicator                           - conditioned for OLLM
    input             PT_phyt_tready_stack,     // Destination Ready                              - conditioned for OLLM
    output [63:0]     BT_phyt_tdata_stack,      // Packet for transfer                            - conditioned for OLLM
    output [7:0]      BT_phyt_tkeep_stack,      // Byte Enable for transferred packet             - conditioned for OLLM
    output            BT_phyt_tlast_stack,      // Last DW of incoming packet                     - conditioned for OLLM
    output [7:0]      BT_phyt_tuser_stack,      // {1'b0, SKIP_CRC, 2'h00, VC[1:0], CRF, SRC_DSC} - conditioned for OLLM
    
    output            PT_phy_rewind,            // rewind indicator
    input             PT_phy_rewind_int         // rewind indicator
    // }}} end Port Declarations
  );                  

  generate if (BYPASS == 1) begin: wirethrough_gen
  // {{{ Wirethrough option
    assign BT_phyt_tvalid_stack = BT_phyt_tvalid;
    assign BT_phyt_tdata_stack  = BT_phyt_tdata;
    assign BT_phyt_tkeep_stack  = BT_phyt_tkeep;
    assign BT_phyt_tlast_stack  = BT_phyt_tlast;
    assign BT_phyt_tuser_stack  = BT_phyt_tuser;

    assign PT_phyt_tready       = PT_phyt_tready_stack;
  assign PT_phy_rewind          = PT_phy_rewind_int;
  // }}} end Wirethrough option

  end else begin: no_wirethrough_gen

  // {{{ Wire Declarations
  
  reg           phy_rst_q;

  wire  [80:0]  data_stage0 = {BT_phyt_tkeep, BT_phyt_tlast, BT_phyt_tuser, BT_phyt_tdata};
  reg   [80:0]  data_stage1;
  reg   [80:0]  data_stage2;
  reg   [80:0]  data_stage3;
  reg   [80:0]  data_stage4;
  reg   [80:0]  data_stage5;

  wire          data_valid_stage0 = PT_phyt_tready && BT_phyt_tvalid;
  reg           data_valid_stage1;
  reg           data_valid_stage2;
  reg           data_valid_stage3;
  reg           data_valid_stage4;
  reg           data_valid_stage5;

  reg           flush_pipe_d, flush_pipe;
  reg           pt_phy_rewind_int_q;
  reg           eop_stack_q;
  reg           allow_ready;
  reg           allow_ready_delay;
  reg           stack_full;
  reg           in_packet;
  reg           in_packet_stack;
  // }}} end Wire Declarations


  // {{{ Register Reset
  // Must register the reset before use
  always @(posedge phy_clk) begin
    phy_rst_q <= #TCQ phy_rst;
  end  
  // }}} end Register Reset


  // {{{ Simple assignments

  assign BT_phyt_tkeep_stack = data_stage5[80:73];
  assign BT_phyt_tlast_stack = data_stage5[72];
  assign BT_phyt_tuser_stack = data_stage5[71:64];
  assign BT_phyt_tdata_stack = data_stage5[63:0];

  assign BT_phyt_tvalid_stack = data_valid_stage5;

  assign PT_phyt_tready = !stack_full;
  assign PT_phy_rewind = PT_phy_rewind_int || allow_ready_delay || allow_ready;
  // }}} end Simple assignments


  // {{{ Flush conditions
  // Clear the pipe after a rewind is observed, but only after tlast gets sent
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      in_packet_stack <= #TCQ 1'b0;
    end else if (BT_phyt_tvalid_stack && !(PT_phyt_tready_stack && BT_phyt_tlast_stack)) begin
      in_packet_stack <= #TCQ 1'b1;
    end else if (BT_phyt_tvalid_stack && PT_phyt_tready_stack && BT_phyt_tlast_stack) begin
      in_packet_stack <= #TCQ 1'b0;
    end
  end
  always @* begin
    if (PT_phy_rewind_int && !pt_phy_rewind_int_q && !(BT_phyt_tvalid_stack || in_packet_stack)) begin
      flush_pipe_d = 1'b1;
    end else if (PT_phy_rewind_int && BT_phyt_tlast_stack && BT_phyt_tvalid_stack && PT_phyt_tready_stack) begin
      flush_pipe_d = 1'b1;
    end else if (PT_phy_rewind_int || allow_ready || allow_ready_delay) begin
      flush_pipe_d = flush_pipe;
    end else begin
      flush_pipe_d = 1'b0;
    end
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      flush_pipe  <= #TCQ 1'b0;
      eop_stack_q <= #TCQ 1'b0;
    end else begin
      flush_pipe  <= #TCQ flush_pipe_d;
      eop_stack_q <= #TCQ BT_phyt_tlast_stack && BT_phyt_tvalid_stack && PT_phyt_tready_stack;
    end
  end



  // }}} end Flush conditions


  // {{{ Valid stages
  wire [5:0] valid_stage = {data_valid_stage5, data_valid_stage4, data_valid_stage3,
                            data_valid_stage2, data_valid_stage1, data_valid_stage0};
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      data_valid_stage5 <= #TCQ 1'b0;
      data_valid_stage4 <= #TCQ 1'b0;
      data_valid_stage3 <= #TCQ 1'b0;
      data_valid_stage2 <= #TCQ 1'b0;
      data_valid_stage1 <= #TCQ 1'b0;
    end else begin
      data_valid_stage5 <= #TCQ ((!PT_phyt_tready_stack && valid_stage[5]) || |valid_stage[4:0]) &&
                                 !(flush_pipe_d || flush_pipe);

      data_valid_stage4 <= #TCQ ((!PT_phyt_tready_stack && valid_stage[4]) ||
                                 (&valid_stage[5:4] && PT_phyt_tready_stack && |valid_stage[3:0]) ||
                                 (valid_stage[5] && !PT_phyt_tready_stack && |valid_stage[3:0])) &&
                                 !flush_pipe;

      data_valid_stage3 <= #TCQ ((!PT_phyt_tready_stack && valid_stage[3]) ||
                                 (&valid_stage[5:3] &&  PT_phyt_tready_stack && |valid_stage[2:0]) ||
                                 (&valid_stage[5:4] && !PT_phyt_tready_stack && |valid_stage[2:0])) &&
                                 !flush_pipe;

      data_valid_stage2 <= #TCQ ((!PT_phyt_tready_stack && valid_stage[2]) ||
                                 (&valid_stage[5:2] &&  PT_phyt_tready_stack && |valid_stage[1:0]) ||
                                 (&valid_stage[5:3] && !PT_phyt_tready_stack && |valid_stage[1:0])) &&
                                 !flush_pipe;

      data_valid_stage1 <= #TCQ ((!PT_phyt_tready_stack && valid_stage[1]) ||
                                 (&valid_stage[5:1] &&  PT_phyt_tready_stack && valid_stage[0]) ||
                                 (&valid_stage[5:2] && !PT_phyt_tready_stack && valid_stage[0])) &&
                                 !flush_pipe;
    end
  end
  // }}} end Valid stages


  // {{{ Data stages
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      data_stage5 <= #TCQ 0;
    end else if (PT_phyt_tready_stack) begin
      casex (valid_stage)
        6'bx1xxxx : data_stage5 <= #TCQ data_stage4;
        default   : data_stage5 <= #TCQ data_stage0;
      endcase
    end else if (!PT_phyt_tready_stack && !valid_stage[5]) begin
      data_stage5 <= #TCQ data_stage0;
    end
  end

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      data_stage4 <= #TCQ 0;
    end else if (PT_phyt_tready_stack) begin
      casex (valid_stage)
        6'bxx1xxx : data_stage4 <= #TCQ data_stage3;
        default   : data_stage4 <= #TCQ data_stage0;
      endcase
    end else if (!PT_phyt_tready_stack && !valid_stage[4]) begin
      data_stage4 <= #TCQ data_stage0;
    end
  end

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      data_stage3 <= #TCQ 0;
    end else if (PT_phyt_tready_stack) begin
      casex (valid_stage)
        6'bxxx1xx : data_stage3 <= #TCQ data_stage2;
        default   : data_stage3 <= #TCQ data_stage0;
      endcase
    end else if (!PT_phyt_tready_stack && !valid_stage[3]) begin
      data_stage3 <= #TCQ data_stage0;
    end
  end

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      data_stage2 <= #TCQ 0;
    end else if (PT_phyt_tready_stack) begin
      casex (valid_stage)
        6'bxxxx1x : data_stage2 <= #TCQ data_stage1;
        default   : data_stage2 <= #TCQ data_stage0;
      endcase
    end else if (!PT_phyt_tready_stack && !valid_stage[2]) begin
      data_stage2 <= #TCQ data_stage0;
    end
  end

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      data_stage1 <= #TCQ 0;
    end else if (PT_phyt_tready_stack) begin
      data_stage1 <= #TCQ data_stage0;
    end else if (!PT_phyt_tready_stack && !valid_stage[1]) begin
      data_stage1 <= #TCQ data_stage0;
    end
  end

  // }}} end Data stages


  // {{{ Full determination

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      pt_phy_rewind_int_q <= #TCQ 1'b0;
    end else begin
      pt_phy_rewind_int_q <= #TCQ PT_phy_rewind_int;
    end
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      in_packet <= #TCQ 1'b0;
    end else if (BT_phyt_tvalid && !(PT_phyt_tready && BT_phyt_tlast)) begin
      in_packet <= #TCQ 1'b1;
    end else if (BT_phyt_tvalid && PT_phyt_tready && BT_phyt_tlast) begin
      in_packet <= #TCQ 1'b0;
    end
  end

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      allow_ready       <= #TCQ 1'b0;
      allow_ready_delay <= #TCQ 1'b0;
    end else if (allow_ready_delay && !valid_stage[3]) begin
      allow_ready       <= #TCQ 1'b1;
      allow_ready_delay <= #TCQ 1'b0;
    end else if (allow_ready && valid_stage[3] && !BT_phyt_tlast) begin
      allow_ready       <= #TCQ 1'b0;
      allow_ready_delay <= #TCQ 1'b1;
    end else if (PT_phy_rewind_int && !pt_phy_rewind_int_q && (BT_phyt_tvalid || in_packet) &&
                 !(BT_phyt_tvalid && PT_phyt_tready && BT_phyt_tlast)) begin
      allow_ready       <= #TCQ !valid_stage[3] || (BT_phyt_tlast && !valid_stage[1]);
      allow_ready_delay <= #TCQ !(!valid_stage[3] || (BT_phyt_tlast && !valid_stage[1]));
    end else if (BT_phyt_tvalid && PT_phyt_tready && BT_phyt_tlast) begin
      allow_ready       <= #TCQ 1'b0;
      allow_ready_delay <= #TCQ 1'b0;
    end
  end


  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      stack_full <= #TCQ 1'b0;
    // create a ready signal that asserts until the last beat of a packet gets through on a rewind
    end else if (allow_ready && !(BT_phyt_tvalid && PT_phyt_tready && BT_phyt_tlast)) begin
      stack_full <= #TCQ 1'b0;
    end else if ((PT_phy_rewind_int || flush_pipe) || allow_ready_delay) begin
      stack_full <= #TCQ 1'b1;
    end else if (&valid_stage[5:1] && !PT_phyt_tready_stack) begin
      stack_full <= #TCQ 1'b1;
    end else if (&valid_stage[5:2] && valid_stage[0] && !PT_phyt_tready_stack) begin
      stack_full <= #TCQ 1'b1;
    end else if (&valid_stage[5:0]) begin
      stack_full <= #TCQ 1'b1;
    end else begin
      stack_full <= #TCQ 1'b0;
    end
  end
  // }}} end Full determination

  end endgenerate

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/phy/ollm_tx/srio_gen2_v4_1_16_ollm_tx_cs_gen.v#1 $
//----------------------------------------------------------------------
//
// OLLM_TX_CS_GEN
// Description:
// This module generates all the control symbols as needed.
//
// Hierarchy:
// PHY_TOP
//    |___OLLM_TX_TOP 
//             |_____OLLM_TX_READY_GEN
//             |_____OLLM_TX_BUF
//             |_____OLLM_TX_PKT_ASSEMBLY
//             |_____OLLM_TX_CS_GEN <-- this module
//             |_____OLLM_TX_DATA_MUX
//             |_____OLLM_TX_OPLM
// ---------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_ollm_tx_cs_gen
  #(
    parameter TCQ         = 100,
    parameter LINK_WIDTH  = 1,    // Generated Link Width {1, 2, 4}
    parameter GT_BYTES    = 4,    // Bytes per cycle on the gt interface
    parameter IDLE1       = 1,    // Include the IDLE1 Sequence {0,1}
    parameter IDLE2       = 0,    // Include the IDLE2 Sequence {0,1}
    parameter VC          = 0,    // Highest numbered VC supported {0,1}
    parameter SIM_TRAIN   = 0)    // {0: FULL, 1: DIVIDED, 3: TRAINED} 
  (
    // {{{ Port Declarations
    // System Signals
    input               phy_clk,                    // PHY interface clock
    input               phy_rst,                    // Reset for PHY clock Domain
    input               log_clk,                    // LOG interface clock
    input               log_rst,                    // Reset for LOG clock Domain
    input               sim_train_en,               // Enable the SIM_TRAIN parameter

    // TX Buffer Interface Signals 
    input               BT_tx_flow_control,         // Indicates the tx buffer is in
                                                    //  tx flow control mode
    
    // RX Buffer Interface Signals
    input       [5:0]   BR_phy_buf_stat,            // VC0 status from the RX buffer 
    input       [5:0]   BR_phy_buf_stat_vc1,        // VC1 status from the RX buffer

    // OPLM TX Interface Signals
    input               PP_port_initialized,        // Indicates port is initialized 
    input               PP_mode_1x,                 // Indicates the link trained down to 1x
    input               PP_idle2_selected,          // Indicated the operating idle mode
    input               PP_ccomp_req,               // Request break for clock comp sequence
    input               PT_ccomp_grant,             // Granted break for clock comp sequence

    // PHY Config Interface Signals
    input               PC_send_lreq,               // Send a Link Request Input Status CS
    input       [2:0]   PC_lreq_cmd,                // Command information for PC_send_lreq
    input               PC_vc_en,                   // Enable VC1
    input       [7:0]   PC_vc1_refresh_int,         // The Refresh Interval for VC1 
    input               PC_load_nextpkt,            // Indicated when a new ackid is loaded in the 
                                                    // ollm rx

    // OLLM RX Interface Signals
    output reg          PTS_sent_init_cs,           // Indicates the link init seq. was sent
    input               PR_send_rfr,                // Send an RFR control symbol 
    output reg          PTS_rfr_sent,               // Sent RFR 
    input               PR_send_lreq,               // Send a Link Request Input Status
    output reg          PTS_lreq_sent,              // Sent Link Request Input Status
    input               PR_send_pna,                // Send a PNA control symbol
    output reg          PTS_pna_sent,               // Sent PNA
    input               PR_send_pr,                 // Send a PR control symbol
    output reg          PTS_pr_sent,                // Sent PR
    input               PR_send_lresp,              // Send a Link Response Control Symbol
    output reg          PTS_lresp_sent,             // Sent Link Response
    
    input       [5:0]   PR_last_good_pkt,           // Last PA to send
    input       [4:0]   PR_cause,                   // Last cause for a PNA to send
    input       [4:0]   PR_port_stat,               // Current port status
    input               PR_link_initialized,        // Link is initialized
    input               PR_output_error_stop,       // Indicates the OLLM RX is in the output error 
                                                    //  stopped state and a LREQ is oustanding
    input               PR_rcvd_error_free_status,  // Indicates when an error free status cs
                                                    // is recieved from the link partner
    // User Interface Signals
    input               UG_phy_mce,                 // Send MCE control symbol 

    // TX Buffer Interface Signals
    input               PTB_in_packet,              // Indicates in packet
    input               PTB_sop,                    // SOP
    input               PTB_eop,                    // EOP
    input               PTB_src_disc,               // source disconnect (mainly for STOMP) // cr 800810, stomp
    input               PTB_sop_d,                  // one cycle early version of PTB_sop
    input       [5:0]   PTB_next_fm,                // The next expected frame's ID
    input               PTR_ptb_advance,            // An active PTB cycle
    input               PTB_link_reset,             // Send link reset control symbols

    // TX Packet Assembly Interface Signals
    input               PTA_in_packet,              // in a packet
    input               PTA_eop,                    // end of a packet
    input       [1:0]   PTA_valid_d,                // Upcoming valid data
    
    // OLLM TX Data Mux Interface 
    output wire [63:0]  PTS_data,                   // Data
    output wire [1:0]   PTS_valid,                  // Valid Data Present on PTS_data
    output wire         PTS_lreq,                   // Indicates the data is a link request
    output wire         PTS_embed_cs,               // Indicates to force the control symbol 
    output wire [7:0]   PTS_charisk,                // Indicates which bytes are K characters 
    output wire         PTS_sop,                    // Indicates the control symbol is an SOP
    output wire         PTS_eop,                    // Indicates the control symbol is an EOP

    // OLLM TX Ready Generator Interface
    output wire         PTS_stall,                  // Stall to PA
    input               PTR_pta_advance,            // Advance the buf interface module
    input               PTR_pts_advance,            // Advance the CS Generator 

    // Output Debug signals
    output reg          PTS_mce_sent,               // Indicates a MCE was sent
    output reg          PTS_pa_sent                 // Indicates a PA was sent
    // }}} end Port Declarations
  );                  

  // {{{ Local Parameters
  // Spec defined parameters
  // ------------------------------------------------------------
  // Stype0
  localparam STYPE0_PA      = 3'b000;
  localparam STYPE0_PR      = 3'b001;
  localparam STYPE0_PNA     = 3'b010;
  localparam STYPE0_STAT    = 3'b100;
  localparam STYPE0_VCSTAT  = 3'b101;
  localparam STYPE0_LRESP   = 3'b110;

  // Stype1
  localparam STYPE1_SOP     = 3'b000;
  localparam STYPE1_STOMP   = 3'b001;// cr 800810, stomp
  localparam STYPE1_EOP     = 3'b010;
  localparam STYPE1_RFR     = 3'b011;
  localparam STYPE1_LREQ    = 3'b100;
  localparam STYPE1_MCE     = 3'b101;
  localparam STYPE1_NOP     = 3'b111;

  //LREQ Commands
  localparam RESET_DEVICE_CMD   = 3'b011;
  localparam INPUT_STATUS_CMD   = 3'b100;
  localparam NO_CMD             = 3'b000;

  // Control Symbol Delimiters
  localparam PD = 8'h7C; //K28.3 8B/10B Character
  localparam SC = 8'h1C; //K28.0 8B/10B Character
 
  // Non-spec. implementation parameters
  // --------------------------------------------------------------
  // The parameter0/1 fields of control symbols are 6-bits in IDLE2
  localparam PARAM_WIDTH  = (IDLE2) ? 6 : 5;

  // The number of outstanding packets you can have in IDLE1 is 32, in IDLE2 its 64
  localparam PA_CTR_WIDTH = (IDLE2) ? 6 : 5;

  // Cycles to space out sending status control symbols for the init sequence
  // Make the timing between the two smaller if the sim_train parameter is set 
  // to divided counters or trained
  // 11 bits is 1024 cycles, 7 bits is 64 cycles
  wire [3:0] INIT_SPACING_WIDTH = (sim_train_en) ? 7 : 11; 

  // Number of outstanding PA's before embedding is required
  localparam EMBED_PA_IDLE1 = 1; // CR 800810 fixed
  localparam EMBED_PA_IDLE2 = 50;

  // Counter length for the codegroups based on the link width
  localparam CG_CTR_WIDTH = (LINK_WIDTH == 4) ? 10 :
                            (LINK_WIDTH == 2) ? 9 : 8;
  localparam CG_TRAINED   = 8;

  // One hot encodings for stype0 functions
  localparam LRESP_ONEHOT             = 6'b10_0000;
  localparam LRESP_BIT                = 5;
  localparam LRESP_BINARY             = 3'h6;

  localparam PNA_ONEHOT               = 6'b01_0000;
  localparam PNA_BIT                  = 4;
  localparam PNA_BINARY               = 3'h5;

  localparam PA_ONEHOT                = 6'b00_1000;  
  localparam PA_BIT                   = 3;  
  localparam PA_BINARY                = 3'h4;

  localparam PR_ONEHOT                = 6'b00_0100;
  localparam PR_BIT                   = 2;
  localparam PR_BINARY                = 3'h3;

  localparam VCSTAT_ONEHOT            = 6'b00_0010;
  localparam VCSTAT_BIT               = 1;
  localparam VCSTAT_BINARY            = 3'h2;

  localparam STAT_ONEHOT              = 6'b00_0001;
  localparam STAT_BIT                 = 0;
  localparam STAT_BINARY              = 3'h1;

  localparam NONE_ONEHOT              = 6'b00_0000;
  localparam NONE_BINARY              = 3'h0;

  // One hot encodings for stype1 functions
  localparam MCE_ONEHOT               = 8'b1000_0000;  
  localparam MCE_BIT                  = 7;  
  localparam MCE_BINARY               = 4'h8;

  localparam CCOMP_EOP_ONEHOT         = 8'b0100_0000;
  localparam CCOMP_EOP_BIT            = 6;
  localparam CCOMP_EOP_BINARY         = 4'h7;

  localparam SOP_ONEHOT               = 8'b0010_0000;
  localparam SOP_BIT                  = 5;
  localparam SOP_BINARY               = 4'h6;

  localparam EOP_ONEHOT               = 8'b0001_0000;
  localparam EOP_BIT                  = 4;
  localparam EOP_BINARY               = 4'h5;

  localparam LREQ_RESET_DEVICE_ONEHOT = 8'b0000_1000;
  localparam LREQ_RESET_DEVICE_BIT    = 3;
  localparam LREQ_RESET_DEVICE_BINARY = 4'h4;

  localparam RFR_ONEHOT               = 8'b0000_0100;
  localparam RFR_BIT                  = 2;
  localparam RFR_BINARY               = 4'h3;

  localparam LREQ_INPUT_STATUS_ONEHOT = 8'b0000_0010;
  localparam LREQ_INPUT_STATUS_BIT    = 1;
  localparam LREQ_INPUT_STATUS_BINARY = 4'h2;

  localparam LREQ_USERDEF_ONEHOT      = 8'b0000_0001;
  localparam LREQ_USERDEF_BIT         = 0;
  localparam LREQ_USERDEF_BINARY      = 4'h1;

  localparam NOP_ONEHOT               = 8'b0000_0000;
  localparam NOP_BINARY               = 4'h0;
  // }}} end Local Parameters
    
  // {{{ Wire Declarations
  reg                     phy_rst_q = 1;
  reg                     log_rst_q = 1;


  // Signals which indicate to send/generate a certain control symbol.
  reg                     send_vcstatus;
  wire                    send_status;
  reg                     send_pa;
  wire                    send_status_init_seq;
  wire                    send_vcstatus_init_seq;
  reg                     send_sop;
  reg                     send_eop;
  wire                    send_lreq;
  wire                    send_rfr;
  reg                     send_ccomp_eop;
  reg                     send_link_reset;
  reg                     link_reset_request;

  //Signals Indicating a sent symbol should be acked.
  wire                    ack_pna;
  wire                    ack_lresp;
  wire                    ack_pr;
  wire                    ack_pa;
  wire                    ack_mce;
  wire                    ack_status;
  wire                    ack_lreq;
  wire                    ack_rfr;
  wire                    ack_eop;

  // Control Symbols Fields for Stype 0 function
  // Default the stype registers in case IDLE2 only and two control symbols 
  // are not being generated.
  reg   [PARAM_WIDTH-1:0] parameter0_0;
  reg   [PARAM_WIDTH-1:0] parameter1_0;
  reg   [PARAM_WIDTH-1:0] parameter0_1;
  reg   [PARAM_WIDTH-1:0] parameter1_1;  
  reg   [2:0]             stype0_0;
  reg   [2:0]             stype0_1;
  reg                     stype0_0_lresp;
  reg                     stype0_0_pa;
  reg                     stype0_0_stat;
  reg                     stype0_0_pna;
  reg                     stype0_0_pr;
  wire  [5:0]             stype0_onehot_0;
  wire  [2:0]             stype0_binary_0;
  wire  [5:0]             stype0_onehot_1;
  reg                     stype0_valid_0;       // Indicates stype0 is valid on the LHS of 64-bit bus
  wire                    stype0_embed;         // Indicates that an stype0 needs to be forced 
  reg                     stype0_embed_q;       // registered stype0_embed 
  wire                    stype0_embed_rose;    // rising edge of stype0_embed 
  reg                     stype0_embed_0;       // Indicates that an stype0 needs to be forced 
  reg   [PARAM_WIDTH-1:0] last_good_pkt_local;  // Local value for current PA param0
  wire                    last_good_pkt_changed;// A change in the last_good_pkt bus
  wire  [PARAM_WIDTH-1:0] param0_last_good_pkt_single;
  wire  [PARAM_WIDTH-1:0] param0_last_good_pkt_multi;
  wire  [PARAM_WIDTH-1:0] param0_last_good_pkt;
  wire  [PARAM_WIDTH-1:0] lresp_last_good_pkt;

  // Control Symbol Fields for an Stype 1 Function
  reg   [2:0]             stype1_0;
  reg   [2:0]             stype1_1;
  reg   [2:0]             stype1_cmd_0;
  reg   [2:0]             stype1_cmd_1;
  reg                     stype1_valid_0;
  reg                     stype1_valid_1;
  wire  [7:0]             stype1_onehot_0;
  wire  [3:0]             stype1_binary_0;
  wire  [7:0]             stype1_onehot_1;
  wire  [3:0]             stype1_binary_1;
  reg                     stype1_embed_0;
  reg                     stype1_embed_1;
  reg                     stype1_0_mce;
  reg                     stype1_eop;
  reg                     stype1_sop;
  reg                     stype1_0_rfr;
  reg                     stype1_0_lreq;
  reg                     stype1_0_lreq_rd;
  reg                     stype1_1_mce;
  reg                     stype1_1_rfr;
  reg                     stype1_1_lreq;
  reg   [7:0]             delimiter_0;
  reg   [7:0]             delimiter_1;

  reg   [4:0]             init_seq_ctr;               // How many init sequence status symbols were sent
  reg                     embed_pa;                   // PAs require embedding
  wire                    buf_stat_int_expired;       // The buf_stat must now be inserted
  reg                     lresp_sent_send_stat;       // Indicates an lresp was sent 
  wire                    assert_send_eop;            // Indicates to end an EOP
  wire                    ending_eop;                 // EOP detected
  wire                    in_packet;                  // A packet is in progress in the OLLM TX
  reg [PA_CTR_WIDTH-1:0]  outstanding_pa_ctr;         // Number of PA to send
  reg                     outstanding_pa_ctr_zero;    //the PA ctr is non-zero
  reg                     outstanding_pa_ctr_one;     //the PA ctr is one
  reg                     send_ccomp_eop_q;           // Registered indicator that a ccomp EOP needs to be sent

  // The control symbol fields to pass to the data mux for
  // both long or short control symbols which are then selected based
  // on the operating idle mode
  wire  [63:0]            short_cs_data;
  wire  [1:0]             short_cs_valid;
  wire                    short_cs_embed;
  wire                    short_cs_lreq;
  wire  [7:0]             short_cs_charisk;
  wire                    short_cs_sop;
  wire                    short_cs_eop;
  reg                     short_cs_stall;
  wire  [63:0]            long_cs_data;
  wire  [1:0]             long_cs_valid;
  wire                    long_cs_embed;  
  wire                    long_cs_lreq;  
  wire  [7:0]             long_cs_charisk;
  wire                    long_cs_sop;
  wire                    long_cs_eop;
  reg                     long_cs_stall;
  // }}} end Wire Declarations

  // {{{ if SIMULATION
  // Make STYPES readable in the waveform for simulation
  `ifdef SIMULATION
    reg [15*8-1:0] stype0_0_string = "null";
    reg [15*8-1:0] stype0_1_string = "null";
    reg [15*8-1:0] stype1_0_string = "null";
    reg [15*8-1:0] stype1_1_string = "null";
    reg [15*8-1:0] cs_symbol_string = "null";

    always @* begin
      //STYPE0 Decode
      case (stype0_0)
        STYPE0_PA:     stype0_0_string = "PA";
        STYPE0_PR:     stype0_0_string = "PR";
        STYPE0_PNA:    stype0_0_string = "PNA";
        STYPE0_STAT:   stype0_0_string = "STAT";
        STYPE0_VCSTAT: stype0_0_string = "VC_STAT";
        STYPE0_LRESP:  stype0_0_string = "LRESP";
        default:       stype0_0_string = "INVALID";
      endcase
      //STYPE1 Decode
      case (stype1_0)
        STYPE1_SOP:  stype1_0_string = "SOP";
        STYPE1_EOP:  stype1_0_string = "EOP";
        STYPE1_RFR:  stype1_0_string = "RFR";
        STYPE1_LREQ: stype1_0_string = "LREQ";
        STYPE1_MCE:  stype1_0_string = "MCE";
        STYPE1_NOP:  stype1_0_string = "NOP";
        default:     stype1_0_string = "INVALID";
      endcase
      case (stype1_1)
        STYPE1_SOP:  stype1_1_string = "SOP";
        STYPE1_EOP:  stype1_1_string = "EOP";
        STYPE1_RFR:  stype1_1_string = "RFR";
        STYPE1_LREQ: stype1_1_string = "LREQ";
        STYPE1_MCE:  stype1_1_string = "MCE";
        STYPE1_NOP:  stype1_1_string = "NOP";
        default:     stype1_1_string = "INVALID";
      endcase
    end
  `endif
  // }}} if SIMULATION

  // {{{ Register Reset
  // Must register the reset before use
  always @(posedge phy_clk) begin
    phy_rst_q <= #TCQ phy_rst;
  end
  always @(posedge log_clk) begin
    log_rst_q <= #TCQ log_rst;
  end
  // }}} end Register Reset

  // {{{ Initialization Sequence
  // Prior to link initialization 15 status control symbols must be sent
  // and 1 VC status symbol if VC1 is enabled. 
  reg [10:0]  init_spacing_ctr;

  // Indicate when to send a status/vcstatus control symbol
  // When VC == 0, 16 Status symbols will be sent, 
  // When VC == 1, 15 Status and 1 VC will be sent
  assign send_status_init_seq   = (!init_seq_ctr[4]) && init_spacing_ctr[INIT_SPACING_WIDTH-1]; 
  // REQ: req_pt_vcstatus_before_link_init
  assign send_vcstatus_init_seq = (!VC) ? 0 :
                                   ((init_seq_ctr == 15) && init_spacing_ctr[INIT_SPACING_WIDTH-1]);
  
  // Reset sending the init sequence if port initialized ever drops
  // wait until one error free status has been recieved to begin counting
  // the control symbols that are sent.  Prior to the OLLM RX recieving an
  // error free status, status symbols will still be sent however just not 
  // counted. These are inserted based on the buf_stat_codegroups counter
  // expiring.
  reg init_seq_enable;

  // REQ: req_pt_status_before_link_init
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      init_seq_enable <= #TCQ 0;
    end else begin
      if (!PP_port_initialized) begin
        init_seq_enable <= #TCQ 0;

      end else if (PR_rcvd_error_free_status) begin
        init_seq_enable <= #TCQ 1'b1;
      end
    end
  end

  // Counter Initialization Sequence Control Symbols Sent
  wire init_seq_ctr_rst     = !init_seq_enable && !PR_rcvd_error_free_status;

  reg advance_init_seq_ctr;

  always @(posedge phy_clk) begin
    advance_init_seq_ctr <= #TCQ !init_seq_ctr[4] && PTR_pts_advance && |PTS_valid;
  end

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      init_seq_ctr <= #TCQ 0;
    end else begin
      // Reset sending the init sequence if port initialized ever drops
      if (init_seq_ctr_rst) begin
        init_seq_ctr <= #TCQ 0;

      // Whenever a control symbol is accepted, increment the counter
      // hold the value when 16
      end else if (advance_init_seq_ctr) begin
        init_seq_ctr <= #TCQ init_seq_ctr + 1'b1;
      end
    end
  end

  //*ASSERTION*
  //(ap_init_seq_ctr_countover): The init_seq_ctr can not count pass 16 

  //*COVERAGE*
  //(cp_init_resets_before_link_init):  Cover that the port_initialized drops
  //before the init_seq_ctr reaches 16.

  //*COVERAGE*
  //(cp_link_init_cycles): Cover that the link initializes from 1-100 cycles after 
  //PTS_sent_init_cs asserts.

  //*ASSERTION*
  //(ap_init_seq_ctr_overcount): The init_seq_ctr can not count past 16

  //*COVERAGE*
  //(cp_vcstatus_during_init): When VC==1, cover that a vc status is sent in init
  //as well as doesn't get sent in init based on PC_vc_en

  // Count based on the init_spacing parameter before sending the next status
  // control symbol.  Reset once the symbol is inserted or port init drops
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      init_spacing_ctr <= #TCQ 0;
    end else begin
      if ((|PTS_valid && PTR_pts_advance) || !PP_port_initialized || !init_seq_enable) begin
        init_spacing_ctr <= #TCQ 0;

      end else if (!init_spacing_ctr[INIT_SPACING_WIDTH-1])begin
        init_spacing_ctr <= #TCQ init_spacing_ctr + 1'b1;
      end
    end
  end
  //*ASSERTION*
  //(ap_init_spacing_ctr_rollsover): The init_spacing_ctr can not roll over.
  
  // We have sent the init sequence as long as the count reaches 16
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PTS_sent_init_cs <= #TCQ 0;
    end else begin
      PTS_sent_init_cs <= #TCQ init_seq_ctr[4];
    end
  end
  // }}} end Initialization Sequence

  // {{{ Stype0 Function Generator
  // The stype0 generator generates stype0 functions with the 
  // following priority:
  // 1. LRESP  (link-response)
  // 2. PNA    (packet-not-accepted)
  // 3. PA     (packet-accepted)
  // 4. PR     (packet-retry)
  // 5. VCSTAT (vc-status)
  // 6. STATUS (status)

  // Only request a send if it wasnt just sent
  wire send_lresp = (PR_send_lresp && !PTS_lresp_sent) && !ack_lresp && !lresp_sent_send_stat;
  
  reg send_pna_d;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      send_pna_d   <= #TCQ 0;
    end else begin

      if (ack_pna || PTS_pna_sent) begin
        send_pna_d <= #TCQ 0;
      end else if (PR_send_pna) begin
        send_pna_d <= #TCQ 1;
      end
    end
  end

  wire send_pna = send_pna_d && !ack_pna;

  // For PR's if a PA is recieved at the same time, we need to wait to send the
  // PA then the PR since there can be no outstanding PAs at the time a PR is
  // sent.
  // Register the PR_send_pr signal so it remains in line with the last_good_pkt_changed signal
  // this helps with timing. 
  reg send_pr_d;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      send_pr_d   <= #TCQ 0;
    end else begin

      if (ack_pr || PTS_pr_sent || last_good_pkt_changed) begin
        send_pr_d <= #TCQ 0;

      end else if (outstanding_pa_ctr_zero && PR_send_pr) begin
        send_pr_d <= #TCQ 1;
      end
    end
  end
  
  wire send_pr = send_pr_d && !ack_pr && !PR_send_pna;

  //*COVERAGE*
  //(cp_pr_and_pna_assert): Cover that PR_send_pr and PR_send_pna assert within various cycles 
  //of eachother 

  //*ASSERTION*
  //(ap_pr_w_outstanding_pna): PR can not assert while there is an outstanding PNA

  // Sort the functions according to their priority left to right
  wire [5:0] stype0_functions_0 = {send_lresp, send_pna, send_pa, 
                                   send_pr, send_vcstatus, send_status};

  //*COVERAGE* 
  //(cr_stype0_functions): Cross all the stype0 functions:
  //PR_send_lresp, PR_send_pna, send_pa, PR_send_pr, send_vcstatus, send_status
  //illegal bins are lresp can never assert with a PNA or a PR
  
  // Get the onehot/binary versions of the function to send
  assign stype0_onehot_0 = stype0_onehot(stype0_functions_0, stype0_embed);
  assign stype0_binary_0 = stype0_binary(stype0_functions_0, stype0_embed);

  // Mask off the buf_stat to all 1's if we are in RX Flow Control
  reg [PARAM_WIDTH-1:0] buf_stat;
  reg [PARAM_WIDTH-1:0] buf_stat_vc1;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      buf_stat     <= #TCQ -1;
      buf_stat_vc1 <= #TCQ -1;
    end else begin
      buf_stat     <= #TCQ (BT_tx_flow_control) ? BR_phy_buf_stat     : -1;
      buf_stat_vc1 <= #TCQ (BT_tx_flow_control) ? BR_phy_buf_stat_vc1 : -1;
    end
  end

  //*COVERAGE*
  //(cp_tx_flow_ctrl): Cover both values of BT_tx_flow_control for sending
  // a PR, PA, STAT or VCSTAT

  //*COVERAGE*
  //(cr_tx_fc_X_idle_selected): Cross the tx flow control signal with PP_idle2_selected.
  
  wire overwrite_pr_pna = (stype0_0 == STYPE0_PR) && (stype0_onehot_0[PNA_BIT]) && 
                          !PTR_pts_advance;

  // Only generate a new symbol if:
  // 1. no symbol is currently valid
  // 2. the valid one has been accepted
  // 3. the special case of a PNA overwritting a PR 
  // 4. the special case of needing to insert an embedded control symbol
  // Nothing should be sent with a LREQ since this could results in multiple
  // cs's going out incorrectly for x1 cores. Mask off stype0 in that case
  // which is ok because the user is trying to bring down the link anyway so
  // that control symbol doesnt need to be sent.
  wire advance_stype0 = (!stype0_valid_0 || PTR_pts_advance || overwrite_pr_pna || stype0_embed_rose) &&
                        !stype1_0_lreq_rd;
 
  // Generate the embed flag with the symbol
  // Need to force the symbol if 
  // 1. the buffer status hasnt been inserted in a while
  // 2. ack ids are running low
  // 3. sending a PNA, all pna's should be embedded for a quick turn
  //    around time.
  // 4. sending a PR, all pr's should be embedded for a quick turn
  //    around time.
  assign stype0_embed = (buf_stat_int_expired && !ack_status) || embed_pa || send_pna || send_pr;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      stype0_embed_q <= #TCQ 0;
    end else begin
      stype0_embed_q <= #TCQ stype0_embed;
    end
  end

  assign stype0_embed_rose = stype0_embed && !stype0_embed_q;

  wire stype0_embed_req_0 = (stype0_onehot_0[STAT_BIT] && buf_stat_int_expired) || 
                            (stype0_onehot_0[PA_BIT]   && embed_pa) ||
                             stype0_onehot_0[PNA_BIT] ||
                             stype0_onehot_0[PR_BIT];

  // Based on the selected stype0, generate the function fields
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      parameter0_0    <= #TCQ 0;
      parameter1_0    <= #TCQ 0;
      stype0_0        <= #TCQ STYPE0_STAT;
      stype0_valid_0  <= #TCQ 0;
      stype0_embed_0  <= #TCQ 0;
      stype0_0_lresp  <= #TCQ 0;
      stype0_0_pa     <= #TCQ 0;
      stype0_0_stat   <= #TCQ 0;
      stype0_0_pna    <= #TCQ 0;
      stype0_0_pr     <= #TCQ 0;

    end else begin
      // Continuously update the CS parameters to have the lateset buf_stat
      // value by the time it is accepted
      // Do not do this for parameter0_1 since it contains acking
      // information which should not get out of sync
      // Do not update if we are not a buf stat (PNAs or LRESPs) and not advancing
      if (advance_stype0) begin
        parameter1_0    <= #TCQ stype0_param1(stype0_binary_0);
      end else if (!stype0_0_pna && !stype0_0_lresp) begin
        parameter1_0    <= #TCQ buf_stat;
      end

      if (advance_stype0) begin
        parameter0_0    <= #TCQ stype0_param0(stype0_binary_0, 
                                              lresp_last_good_pkt, param0_last_good_pkt, PTB_next_fm);
        stype0_0        <= #TCQ stype0_type(stype0_binary_0);
        stype0_valid_0  <= #TCQ |stype0_onehot_0;
        stype0_embed_0  <= #TCQ stype0_embed_req_0;

        // Save off the type of control symbol to improve timing
        stype0_0_lresp  <= #TCQ stype0_onehot_0[LRESP_BIT];
        stype0_0_pa     <= #TCQ stype0_onehot_0[PA_BIT];
        stype0_0_stat   <= #TCQ stype0_onehot_0[STAT_BIT] || ~(|stype0_onehot_0);
        stype0_0_pna    <= #TCQ stype0_onehot_0[PNA_BIT];
        stype0_0_pr     <= #TCQ stype0_onehot_0[PR_BIT];

      end
    end
  end

  //*ASSERTION*
  //(ap_buf_stat5_invalid): if we are in idle1 mode BR_phy_buf_stat[5] must always be 0
  
  //*ASSERTION*
  //(ap_buf_statvc15_invalid): if we are in idle1 mode BR_phy_buf_stat_vc1[5] must always be 0
    always @(posedge phy_clk) begin
      parameter0_1    <= #TCQ PTB_next_fm[PARAM_WIDTH-1:0];
      parameter1_1    <= #TCQ buf_stat;
      stype0_1        <= #TCQ STYPE0_STAT;
    end    

  //*ASSERTION*
  //(ap_rogue_stype0_embed_0): stype0_embed_0 can not assert with no valid control symbols

  // In TX flow control mode an lresp must be followed by a vc status and
  // a status control symbol in that order.  Only ask the lresp after the
  // entire sequence is sent in this mode.
  assign ack_lresp  = (stype0_0_lresp) && PTR_pts_advance;
  
  //Need to be sure that status was valid since this is the filler control
  //symbol
  assign ack_status = (stype1_valid_1 || 
                       (stype0_0_stat && (stype0_valid_0 || stype1_valid_0))) && 
                      PTR_pts_advance;
  
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      lresp_sent_send_stat <= #TCQ 0;
    end else begin
      if (ack_status) begin
        lresp_sent_send_stat <= #TCQ 0;
      end else if (ack_lresp && BT_tx_flow_control) begin
        lresp_sent_send_stat <= #TCQ 1;
      end
    end
  end

  // Acknowledge control symbol requests if they were requested by the OLLM RX
  assign ack_pna = stype0_0_pna && PTR_pts_advance;

  // A PR needs to be acked when a PNA replaces it
  assign ack_pr  = (stype0_0_pr && PTR_pts_advance) ||
                   (ack_pna && PR_send_pr && !PTS_pr_sent);

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PTS_pna_sent   <= #TCQ 0;
      PTS_pr_sent    <= #TCQ 0;
      PTS_lresp_sent <= #TCQ 0;
    end else begin
      PTS_pna_sent   <= #TCQ ack_pna;
      PTS_pr_sent    <= #TCQ ack_pr;
      PTS_lresp_sent <= #TCQ ack_lresp;     
    end
  end 
   
  //*COVERAGE*
  //(cp_pna_overwrites_pr): Cover that a PNA overwrites a PR

  //*ASSERTION*
  //(ap_pna_and_pr_both_acked): When a PNA overwrite a PR both should be acked.

  // {{{ + STYPE0 Utility Functions +
  // {{{ stype0_type -
  // returns the stype field given the one hot encoding
  // REQ: req_pt_buf_stat_sent_as_needed
  function [2:0] stype0_type (
    input [2:0] functions
  ); begin
      case (functions)
        LRESP_BINARY:  stype0_type = STYPE0_LRESP;
        PNA_BINARY:    stype0_type = STYPE0_PNA;
        PA_BINARY:     stype0_type = STYPE0_PA;
        PR_BINARY:     stype0_type = STYPE0_PR;
        VCSTAT_BINARY: stype0_type = STYPE0_VCSTAT;
        STAT_BINARY:   stype0_type = STYPE0_STAT;
        NONE_BINARY:   stype0_type = STYPE0_STAT;
        default:       stype0_type = {3{1'bX}};
      endcase
    end
  endfunction
  // }}} end stype0_type

  // {{{ stype0_param0 -
  // returns the parameter0 field given the one hot encoding

  // If we are using the last good packet in parameter 0, then we need to
  // manage the rollover case for IDLE1 mode.
  assign param0_last_good_pkt_single = (!PP_idle2_selected && (last_good_pkt_local == 31)) ? 0 : 
                                                                                             last_good_pkt_local + 1;

  assign param0_last_good_pkt_multi = (!PP_idle2_selected && (last_good_pkt_local == 31)) ? 1 : 
                                      (!PP_idle2_selected && (last_good_pkt_local == 30)) ? 0 : 
                                                                                            last_good_pkt_local + 2;

  assign param0_last_good_pkt = (ack_pa) ? param0_last_good_pkt_multi : 
                                           param0_last_good_pkt_single;

  assign lresp_last_good_pkt = (!PP_idle2_selected && (PR_last_good_pkt == 31)) ? 0 : 
                                                                                  PR_last_good_pkt + 1;

  function [PARAM_WIDTH-1:0] stype0_param0 (
    input [2:0]             functions,
    input [PARAM_WIDTH-1:0] lresp_last_good_pkt,
    input [PARAM_WIDTH-1:0] param0_last_good_pkt,
    input [5:0]             PTB_next_fm 
  ); begin
      //Only grab the appropriate width for this configuration
      //to avoid truncation warnings in XST.
      case (functions)
        LRESP_BINARY:  stype0_param0 = lresp_last_good_pkt[PARAM_WIDTH-1:0]; 
        PNA_BINARY:    stype0_param0 = {PARAM_WIDTH{1'b0}};
        PA_BINARY:     stype0_param0 = param0_last_good_pkt[PARAM_WIDTH-1:0];
        PR_BINARY:     stype0_param0 = param0_last_good_pkt[PARAM_WIDTH-1:0];
        VCSTAT_BINARY: stype0_param0 = {PARAM_WIDTH{1'b0}};
        //STAT_BINARY:   stype0_param0 = PTB_next_fm[PARAM_WIDTH-1:0];      // this was original logic, CR # 764307 
	    STAT_BINARY:   stype0_param0 = lresp_last_good_pkt[PARAM_WIDTH-1:0];// this is updated to fix the CR # 764307 
        //  NONE_BINARY:   stype0_param0 = PTB_next_fm[PARAM_WIDTH-1:0];
        NONE_BINARY:   stype0_param0 = lresp_last_good_pkt[PARAM_WIDTH-1:0]; // fix for CR # 764307
        default:       stype0_param0 = {PARAM_WIDTH{1'bX}};
      endcase
    end
  endfunction
  // }}} end stype0_param0

  // {{{ stype0_param1 -
  // returns the parameter1 field given the one hot encoding
  function [PARAM_WIDTH-1:0] stype0_param1 (
    input [2:0] functions
  ); begin
      case (functions)
        LRESP_BINARY:  stype0_param1 = {1'b0, PR_port_stat};
        PNA_BINARY:    stype0_param1 = {1'b0, PR_cause};
        PA_BINARY:     stype0_param1 = buf_stat;
        PR_BINARY:     stype0_param1 = buf_stat;
        VCSTAT_BINARY: stype0_param1 = buf_stat_vc1;
        STAT_BINARY:   stype0_param1 = buf_stat;
        NONE_BINARY:   stype0_param1 = buf_stat;
        default:       stype0_param1 = {PARAM_WIDTH{1'bX}};
      endcase
    end
  endfunction
  // }}} end stype0_param1  

  // {{{ stype0_onehot -
  // returns the one hot encoding of the valid stype0 functions
  function [5:0] stype0_onehot (
    input [5:0] functions,
    input       stype0_embed
  ); begin
      casex ({stype0_embed, functions})
        // original code before CR# 725569, // 1/12/2015
	// {1'b0, 6'b1x_xxxx}: stype0_onehot = LRESP_ONEHOT;
        // {1'b1, 6'b01_xxxx}: stype0_onehot = PNA_ONEHOT;
        // {1'b0, 6'b00_1xxx}: stype0_onehot = PA_ONEHOT;   
        // {1'b1, 6'bxx_1xxx}: stype0_onehot = PA_ONEHOT;//it was 6'bxx_1xxx, CR #725569
        // {1'b1, 6'b00_01xx}: stype0_onehot = PR_ONEHOT;
        // {1'b0, 6'b00_001x}: stype0_onehot = VCSTAT_ONEHOT;
        // {1'b0, 6'b00_0001}: stype0_onehot = STAT_ONEHOT;
        // {1'b1, 6'bxx_0xx1}: stype0_onehot = STAT_ONEHOT;// it was 6'bxx_0xx1, CR #725569
        // default           : stype0_onehot = NONE_ONEHOT;

	//****************************************
        // below is the updated code to fix the issue observed in CR# 725569, // 1/12/2015
	{1'b0, 6'b1x_xxxx}: stype0_onehot = LRESP_ONEHOT;
      //{1'b1, 6'b01_xxxx}: stype0_onehot = PNA_ONEHOT;
        {1'b1, 6'b01_0000}: stype0_onehot = PNA_ONEHOT;
        {1'b1, 6'b01_0001}: stype0_onehot = PNA_ONEHOT;
        {1'b1, 6'b01_0010}: stype0_onehot = PNA_ONEHOT;
        {1'b1, 6'b01_0011}: stype0_onehot = PNA_ONEHOT;
        {1'b1, 6'b01_0100}: stype0_onehot = PNA_ONEHOT;
        {1'b1, 6'b01_0101}: stype0_onehot = PNA_ONEHOT;
        {1'b1, 6'b01_0110}: stype0_onehot = PNA_ONEHOT;
        {1'b1, 6'b01_0111}: stype0_onehot = PNA_ONEHOT;
      // {1'b1, 6'b01_1000}: stype0_onehot = PNA_ONEHOT;
      // {1'b1, 6'b01_1001}: stype0_onehot = PNA_ONEHOT;
      // {1'b1, 6'b01_1010}: stype0_onehot = PNA_ONEHOT;
      // {1'b1, 6'b01_1011}: stype0_onehot = PNA_ONEHOT;
      // {1'b1, 6'b01_1100}: stype0_onehot = PNA_ONEHOT;
      // {1'b1, 6'b01_1101}: stype0_onehot = PNA_ONEHOT;
      // {1'b1, 6'b01_1110}: stype0_onehot = PNA_ONEHOT;
      // {1'b1, 6'b01_1111}: stype0_onehot = PNA_ONEHOT;
        {1'b0, 6'b00_1xxx}: stype0_onehot = PA_ONEHOT;   

      //{1'b1, 6'bxx_1xxx}: stype0_onehot = PA_ONEHOT;//it was 6'bxx_1xxx, CR #725569
        {1'b1, 6'b00_1000}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b00_1001}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b00_1010}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b00_1011}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b00_1100}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b00_1101}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b00_1110}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b00_1111}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b01_1000}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b01_1001}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b01_1010}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b01_1011}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b01_1100}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b01_1101}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b01_1110}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b01_1111}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b10_1000}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b10_1001}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b10_1010}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b10_1011}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b10_1100}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b10_1101}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b10_1110}: stype0_onehot = PA_ONEHOT;
        {1'b1, 6'b10_1111}: stype0_onehot = PA_ONEHOT;

      //{1'b1, 6'b00_01xx}: stype0_onehot = PR_ONEHOT;
        {1'b1, 6'b00_0100}: stype0_onehot = PR_ONEHOT;
      //{1'b1, 6'b00_0101}: stype0_onehot = PR_ONEHOT;
        {1'b1, 6'b00_0110}: stype0_onehot = PR_ONEHOT;
      //{1'b1, 6'b00_0111}: stype0_onehot = PR_ONEHOT;

        {1'b0, 6'b00_001x}: stype0_onehot = VCSTAT_ONEHOT;
        {1'b0, 6'b00_0001}: stype0_onehot = STAT_ONEHOT;
        
      //{1'b1, 6'bxx_0xx1}: stype0_onehot = STAT_ONEHOT;// it was 6'bxx_0xx1, CR #725569
	{1'b1, 6'b00_0001}: stype0_onehot = STAT_ONEHOT;// it was 6'bxx_0xx1, CR #725569
	{1'b1, 6'b00_0011}: stype0_onehot = STAT_ONEHOT;// it was 6'bxx_0xx1, CR #725569
	{1'b1, 6'b00_0101}: stype0_onehot = STAT_ONEHOT;// it was 6'bxx_0xx1, CR #725569
	{1'b1, 6'b00_0111}: stype0_onehot = STAT_ONEHOT;// it was 6'bxx_0xx1, CR #725569

	//{1'b1, 6'b01_0001}: stype0_onehot = STAT_ONEHOT;// it was 6'bxx_0xx1, CR #725569
	//{1'b1, 6'b01_0011}: stype0_onehot = STAT_ONEHOT;// it was 6'bxx_0xx1, CR #725569
	//{1'b1, 6'b01_0101}: stype0_onehot = STAT_ONEHOT;// it was 6'bxx_0xx1, CR #725569
	//{1'b1, 6'b01_0111}: stype0_onehot = STAT_ONEHOT;// it was 6'bxx_0xx1, CR #725569

	{1'b1, 6'b10_0001}: stype0_onehot = STAT_ONEHOT;// it was 6'bxx_0xx1, CR #725569
	{1'b1, 6'b10_0011}: stype0_onehot = STAT_ONEHOT;// it was 6'bxx_0xx1, CR #725569
	{1'b1, 6'b10_0101}: stype0_onehot = STAT_ONEHOT;// it was 6'bxx_0xx1, CR #725569
	{1'b1, 6'b10_0111}: stype0_onehot = STAT_ONEHOT;// it was 6'bxx_0xx1, CR #725569

	{1'b1, 6'b11_0001}: stype0_onehot = STAT_ONEHOT;// it was 6'bxx_0xx1, CR #725569
	{1'b1, 6'b11_0011}: stype0_onehot = STAT_ONEHOT;// it was 6'bxx_0xx1, CR #725569
	{1'b1, 6'b11_0101}: stype0_onehot = STAT_ONEHOT;// it was 6'bxx_0xx1, CR #725569
	{1'b1, 6'b11_0111}: stype0_onehot = STAT_ONEHOT;// it was 6'bxx_0xx1, CR #725569

        default           : stype0_onehot = NONE_ONEHOT;
	//****************************************
      endcase
    end 
  endfunction
  // }}} end stype0_onehot

  // {{{ stype0_binary -
  // returns the one hot encoding of the valid stype0 functions
  function [2:0] stype0_binary (
    input [5:0] functions,
    input       stype0_embed
  ); begin
      // If a status needs to be embedded it take priority over any other
      // stype 0 which needs embedding.
      casex ({stype0_embed, functions})
        // original code before CR# 725569, // 1/12/2015
        // {1'b0, 6'b1x_xxxx}: stype0_binary = LRESP_BINARY;
        // {1'b1, 6'b01_xxxx}: stype0_binary = PNA_BINARY;
        // {1'b0, 6'b00_1xxx}: stype0_binary = PA_BINARY;   
        // {1'b1, 6'bxx_1xxx}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        // {1'b1, 6'b00_01xx}: stype0_binary = PR_BINARY;
        // {1'b0, 6'b00_001x}: stype0_binary = VCSTAT_BINARY;
        // {1'b0, 6'b00_0001}: stype0_binary = STAT_BINARY;
        // {1'b1, 6'bxx_0xx1}: stype0_binary = STAT_BINARY;//it was 6'bxx_0xx1 , CR #725569
        // default           : stype0_binary = NONE_BINARY;
      //*******************
        // below is the updated code to fix the issue observed in CR# 725569, // 1/12/2015
        {1'b0, 6'b1x_xxxx}: stype0_binary = LRESP_BINARY;
      //{1'b1, 6'b01_xxxx}: stype0_binary = PNA_BINARY;
        {1'b1, 6'b01_0000}: stype0_binary = PNA_BINARY;
        {1'b1, 6'b01_0001}: stype0_binary = PNA_BINARY;
        {1'b1, 6'b01_0010}: stype0_binary = PNA_BINARY;
        {1'b1, 6'b01_0011}: stype0_binary = PNA_BINARY;
        {1'b1, 6'b01_0100}: stype0_binary = PNA_BINARY;
        {1'b1, 6'b01_0101}: stype0_binary = PNA_BINARY;
        {1'b1, 6'b01_0110}: stype0_binary = PNA_BINARY;
        {1'b1, 6'b01_0111}: stype0_binary = PNA_BINARY;
      //{1'b1, 6'b01_1000}: stype0_binary = PNA_BINARY;
      //{1'b1, 6'b01_1001}: stype0_binary = PNA_BINARY;
      //{1'b1, 6'b01_1010}: stype0_binary = PNA_BINARY;
      //{1'b1, 6'b01_1011}: stype0_binary = PNA_BINARY;
      //{1'b1, 6'b01_1100}: stype0_binary = PNA_BINARY;
      //{1'b1, 6'b01_1101}: stype0_binary = PNA_BINARY;
      //{1'b1, 6'b01_1110}: stype0_binary = PNA_BINARY;
      //{1'b1, 6'b01_1111}: stype0_binary = PNA_BINARY;

        {1'b0, 6'b00_1xxx}: stype0_binary = PA_BINARY;   
      //{1'b1, 6'bxx_1xxx}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b00_1000}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b00_1001}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b00_1010}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b00_1011}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b00_1100}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b00_1101}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b00_1110}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b00_1111}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569

        {1'b1, 6'b01_1000}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b01_1001}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b01_1010}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b01_1011}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b01_1100}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b01_1101}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b01_1110}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b01_1111}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569

        {1'b1, 6'b10_1000}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b10_1001}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b10_1010}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b10_1011}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b10_1100}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b10_1101}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b10_1110}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b10_1111}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569

	{1'b1, 6'b11_1000}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b11_1001}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b11_1010}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b11_1011}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b11_1100}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b11_1101}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b11_1110}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569
        {1'b1, 6'b11_1111}: stype0_binary = PA_BINARY;//it was 6'bxx_1xxx , CR #725569

        //{1'b1, 6'b00_01xx}: stype0_binary = PR_BINARY;
	{1'b1, 6'b00_0100}: stype0_binary = PR_BINARY;
      //{1'b1, 6'b00_0101}: stype0_binary = PR_BINARY;
	{1'b1, 6'b00_0110}: stype0_binary = PR_BINARY;
      //{1'b1, 6'b00_0111}: stype0_binary = PR_BINARY;

        {1'b0, 6'b00_001x}: stype0_binary = VCSTAT_BINARY;
        {1'b0, 6'b00_0001}: stype0_binary = STAT_BINARY;

      //{1'b1, 6'bxx_0xx1}: stype0_binary = STAT_BINARY;//it was 6'bxx_0xx1 , CR #725569
        {1'b1, 6'b00_0001}: stype0_binary = STAT_BINARY;//it was 6'bxx_0xx1 , CR #725569
	{1'b1, 6'b00_0011}: stype0_binary = STAT_BINARY;//it was 6'bxx_0xx1 , CR #725569
	{1'b1, 6'b00_0101}: stype0_binary = STAT_BINARY;//it was 6'bxx_0xx1 , CR #725569
	{1'b1, 6'b00_0111}: stype0_binary = STAT_BINARY;//it was 6'bxx_0xx1 , CR #725569

        //{1'b1, 6'b01_0001}: stype0_binary = STAT_BINARY;//it was 6'bxx_0xx1 , CR #725569
	//{1'b1, 6'b01_0011}: stype0_binary = STAT_BINARY;//it was 6'bxx_0xx1 , CR #725569
	//{1'b1, 6'b01_0101}: stype0_binary = STAT_BINARY;//it was 6'bxx_0xx1 , CR #725569
	//{1'b1, 6'b01_0111}: stype0_binary = STAT_BINARY;//it was 6'bxx_0xx1 , CR #725569

        {1'b1, 6'b10_0001}: stype0_binary = STAT_BINARY;//it was 6'bxx_0xx1 , CR #725569
	{1'b1, 6'b10_0011}: stype0_binary = STAT_BINARY;//it was 6'bxx_0xx1 , CR #725569
	{1'b1, 6'b10_0101}: stype0_binary = STAT_BINARY;//it was 6'bxx_0xx1 , CR #725569
	{1'b1, 6'b10_0111}: stype0_binary = STAT_BINARY;//it was 6'bxx_0xx1 , CR #725569

        {1'b1, 6'b11_0001}: stype0_binary = STAT_BINARY;//it was 6'bxx_0xx1 , CR #725569
	{1'b1, 6'b11_0011}: stype0_binary = STAT_BINARY;//it was 6'bxx_0xx1 , CR #725569
	{1'b1, 6'b11_0101}: stype0_binary = STAT_BINARY;//it was 6'bxx_0xx1 , CR #725569
	{1'b1, 6'b11_0111}: stype0_binary = STAT_BINARY;//it was 6'bxx_0xx1 , CR #725569

        default           : stype0_binary = NONE_BINARY;
      //*******************

      
      endcase
    end 
  endfunction
  // }}} end stype0_binary

  // }}} + end STYPE0 Utility Functions +
  
  // }}} end Stype0 Function Generator

  // {{{ PA Generator
  // A PA needs to be sent for every packet that is acked, indicated
  // by a change in PR_last_good_pkt.  When too many PAs are outstanding
  // the symbol must be sent in order to free up Ack IDs in the link partner
  reg [5:0]              last_good_pkt_q;

  assign ack_pa = stype0_0_pa && PTR_pts_advance;
  
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PTS_pa_sent <= #TCQ 0;
    end else begin
      PTS_pa_sent <= #TCQ ack_pa;
    end
  end

  // Monitor last_good_pkt for changes
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      last_good_pkt_q <= #TCQ (IDLE2) ? 6'h3F : 6'h1F; 
    end else begin
      last_good_pkt_q <= #TCQ PR_last_good_pkt;
    end
  end

  // Register PC_load_nextpkt to know when last good pkt changing is actually
  // valid
  reg load_nextpkt_q;
  reg idle2_selected_q;
  reg idle2_mode_changed;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      load_nextpkt_q      <= #TCQ 0;
      idle2_selected_q    <= #TCQ 0;
      idle2_mode_changed  <= #TCQ 0;
    end else begin
      load_nextpkt_q      <= #TCQ PC_load_nextpkt;
      idle2_selected_q    <= #TCQ PP_idle2_selected;
      idle2_mode_changed  <= #TCQ idle2_selected_q != PP_idle2_selected;

    end
  end

  // If a load ACK ids caused a change in last good pkt, then this does not
  // mean send a PA. in this case gate off the last_good_pkt_changed indicator
  assign last_good_pkt_changed = (last_good_pkt_q != PR_last_good_pkt) && !load_nextpkt_q && 
                                 !idle2_mode_changed;


// Generate a pulse to clear outstanding PA count when lresp is triggered. 
// This will allow if PAs to be sent if any packet comes after LREQ and before LRESP is sent
  reg      stype0_0_lresp_delay;
  always @(posedge phy_clk) begin
    if (phy_rst_q) 
       stype0_0_lresp_delay      <= #TCQ 0;
    else 
       stype0_0_lresp_delay      <= #TCQ stype0_0_lresp;
    end


wire stype0_0_lresp_pulse = stype0_0_lresp & !stype0_0_lresp_delay;




  // Counter to see how many times a packet has been accepted.
  // If the number of oustanding packets exceeds the parameters
  // EMBED_PA_IDLE1/EMBED_PA_IDLE2 then it should be embedded
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      outstanding_pa_ctr      <= #TCQ 0;
      outstanding_pa_ctr_zero <= #TCQ 1;
      outstanding_pa_ctr_one  <= #TCQ 0;
    end else begin
      // On an implicit ack condition reset the oustanding counter
      // Implicitly ack on a PNA since an LRESP has to follow a PNA
      // and it will do the implicit acking for us. However it needs to 
      // be cleared before the lresp is sent so that PNAs are not sent
      // while the link partner is in input error and ignoring those PAs
      //
      // Gate sending any PA before link init in case last good pkt changes 
      // because of the idle mode changing from 2 to 1
      if (stype0_0_lresp_pulse || ack_pna) begin
        outstanding_pa_ctr      <= #TCQ 0;
        outstanding_pa_ctr_zero <= #TCQ 1;
        outstanding_pa_ctr_one  <= #TCQ 0;
      end else begin

        //Dont change stage for both an incr/decr condition
        if (ack_pa && last_good_pkt_changed) begin
          outstanding_pa_ctr      <= #TCQ outstanding_pa_ctr;
          outstanding_pa_ctr_zero <= #TCQ outstanding_pa_ctr_zero;
          outstanding_pa_ctr_one  <= #TCQ outstanding_pa_ctr_one;
        // Decrement the counter for every PA sent
        end else if (ack_pa) begin
          outstanding_pa_ctr      <= #TCQ outstanding_pa_ctr - 1'b1;
          outstanding_pa_ctr_zero <= #TCQ (outstanding_pa_ctr == 1);
          outstanding_pa_ctr_one  <= #TCQ (outstanding_pa_ctr == 2);
        // Increment the counter for every good packet seen
        end else if (last_good_pkt_changed) begin
          outstanding_pa_ctr      <= #TCQ outstanding_pa_ctr + 1'b1;
          outstanding_pa_ctr_zero <= #TCQ 0;
          outstanding_pa_ctr_one  <= #TCQ (outstanding_pa_ctr == 0);
        end
      end
    end
  end  

  // Maintain a local count for the last good packet value to use as param0
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      last_good_pkt_local  <= #TCQ -1;

    end else begin
      // On an implicit ack condition update to the most recent last good pkt
      // If a PNA is sent then update this to the pna value,
      if (ack_lresp || ack_pna) begin
        last_good_pkt_local  <= #TCQ PR_last_good_pkt;

      // Whenever a packet is acked, need to update the local last good pkt
      end else if (ack_pa) begin
        last_good_pkt_local <= #TCQ (!PP_idle2_selected && (last_good_pkt_local == 31)) ?
                                    0 : last_good_pkt_local + 1;
      end 
    end
  end   

  //*COVERAGE*
  //(cp_outstanding_pa_ctr_neutral): Cover that PTR_pts_advance, ack_pa, and last_good_pkt_changed
  //are all asserted 

  //*ASSERTION*
  //(ap_outstanding_pa_ctr_neutral): When PTR_pts_advance, ack_pa, and last_good_pkt_changed are
  //all asserted, the counter should not change

  //*ASSERTION*
  //(ap_pa_ctr_overcount_idle1): the PA_ctr does not count past its max value for idle1 mode (31)

  //*ASSERTION*
  //(ap_pa_ctr_overcount_idle2): the PA_ctr does not count past its max value for idle2 mode (63)
  
  //*ASSERTION*
  //(ap_pa_ctr_rollunder): the PA_ctr does not roll under
  
  //*ASSERTION*
  //(ap_pa_ctr_rollover_idle1): the PA_ctr does not roll over in idle1

  //*ASSERTION*
  //(ap_pa_ctr_rollover_idle2): the PA_ctr does not roll over in idle2
  
  //*COVERAGE*
  //(cp_pa_ctr_values): Cover all the values of the oustanding PA's counter

  //*COVERAGE*
  //(cp_implicit_acks): See a couple of implicit ack conditions
  
  // Indicate when to send a PA and if it should be embeddeda PA should not be 
  // sent if the lresp sequence is not being sent. This is because and lresp 
  // must be followed by a vcstatus and status control symbol and the priority 
  // of a PA would interfer with this sequence.  
  // Do not send any PA's if a PNA needs to be sent, a PNA clears all
  // outstanding PA's anyway
  always @* begin
    if ((outstanding_pa_ctr_one && ack_pa) || stype0_0_lresp_pulse  || 
        PR_send_pna || send_link_reset) begin
      send_pa = 0;
    end else begin
      send_pa = !outstanding_pa_ctr_zero && PR_link_initialized;
    end
  end 

  //*COVERAGE*
  //(cp_link_drops_w_outstanding_pa): See link init drop where there are still
  //outstanding PAs to send

  //*ASSERTION*
  //(ap_pa_sent_before_link_init): A PA can not be sent before link init is
  //asserted.
  //
  //*COVERAGE*
  //(ap_lresp_tx_fc): Cover that an lresp needs to be sent in TX Flow control
  
  //*COVERAGE*
  //(cp_lresp_rx_fc): Cover that an lresp needs to be sent in RX Flow control

  //*ASSERTION*
  //(ap_force_pa_sent): If the pa_ctr is greater than EMBED_PA_IDLE1/EMBED_PA_IDLE2
  //a pa must be embedded and embed_pa assert with send_pa.

  //*COVERAGE*
  //(cp_force_pa_sent): A PA is forced to be sent (embedded)

  // Force PA's to be embeded if:
  // 1. they are starting to build up and IDs available could potentially run out. 
  // 2. Also embed if a PR needs to be sent so that we can send the PR as quickly as possible.
  // 3. If the buf status needs to be inserted immediately and we can insert
  //    it by using the PA
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      embed_pa <= #TCQ 0;
    end else begin
      embed_pa <= #TCQ (PP_idle2_selected) ? 
                        (send_pa && ((outstanding_pa_ctr > EMBED_PA_IDLE2) || PR_send_pr ||
                         buf_stat_int_expired)) :
                        (send_pa && ((outstanding_pa_ctr > EMBED_PA_IDLE1) || PR_send_pr || 
                         buf_stat_int_expired));
    end
  end
  // }}} end PA Generator

  // {{{ VC Status Generator
  // Send the vc status symbol if:
  // 1. the init_seq_ctr indicates to by a value of 15
  // 2. the VC counter expires
  // Only generated VC1 logic if VC is set to 1
  generate if (VC == 1) begin: vc_status_gen
    wire                      buf_stat_vc1_changed;
    reg   [5:0]               buf_stat_vc1_q;
    wire                      vc1_refresh_int_expired;
    reg   [CG_CTR_WIDTH-1:0]  vc1_codegroups_ctr;
    reg   [7:0]               vc1_refresh_int_ctr;
    
    // Monitor VC1 for changes to know when to send this symbol
    // REQ: req_pt_vc_stat_changed_and_sent
    assign buf_stat_vc1_changed = (buf_stat_vc1_q != BR_phy_buf_stat_vc1);

    always @(posedge phy_clk) begin
      if (phy_rst_q) begin
        buf_stat_vc1_q <= #TCQ 0;
      end else begin
        buf_stat_vc1_q <= #TCQ BR_phy_buf_stat_vc1;
      end
    end

    wire vc1_trained_max = PP_mode_1x && vc1_codegroups_ctr[CG_TRAINED-1];

    // The Codegroups counter determines how many codegroups have been sent for
    // this link width. A VC Status must be sent every 1024-codegroups.
    // REQ: req_pt_vc_stat_sent_as_needed
    always @(posedge phy_clk) begin
      if (phy_rst_q) begin
        vc1_codegroups_ctr <= #TCQ 0;
      end else begin
        // When trained, reduce the max count value
        if (vc1_trained_max) begin
          vc1_codegroups_ctr <= #TCQ 0;
        end else begin
          vc1_codegroups_ctr <= #TCQ vc1_codegroups_ctr + 1'b1;
        end
      end
    end

    // Count up until the refresh interval before sending a vc_status
    // this is the multiplier of the codegroup counter.
    always @(posedge phy_clk) begin
      if (phy_rst_q) begin
        vc1_refresh_int_ctr <= #TCQ 0;
      end else begin
        if (vc1_codegroups_ctr[CG_CTR_WIDTH-1] || vc1_trained_max) begin
          vc1_refresh_int_ctr <= #TCQ  + 1'b1;
        end
      end
    end

    // Indicate to send the a VC status if:
    // 1. the send refresh timer timesout
    // 2. the init sequence indicated to send one
    // 2. the buf status for VC1 changes
    // 3. AND PC_vc_en is true.
    // REQ: req_pt_vc_refresh_int_valid
    assign vc1_refresh_int_expired = (vc1_refresh_int_ctr == PC_vc1_refresh_int);
    wire   assert_send_vcstatus    = (send_vcstatus_init_seq || buf_stat_vc1_changed || 
                                      vc1_refresh_int_expired) && PC_vc_en;
    wire   ack_vcstatus            = ((stype0_1 == STYPE0_VCSTAT) || 
                                      (stype0_0 == STYPE0_VCSTAT)) && PTR_pts_advance;

    always @(posedge phy_clk) begin
      if (phy_rst_q) begin
        send_vcstatus <= #TCQ 0;
      end else begin
        // Reset once it is sent
        if (ack_vcstatus) begin
          send_vcstatus <= #TCQ 0;
        end else if (assert_send_vcstatus)  begin
          send_vcstatus <= #TCQ 1;
        end
      end
    end

    //*COVERAGE*
    //(cp_vc1_cg_ctr_expires): A VC status symbol needs to be sent by the
    //timer expiring (vc1_refresh_int_expired).
  
  // When only VC0 is supported tie off sending a vcstatus
  end else begin: no_vc_status_gen
    always @(posedge phy_clk) begin
      send_vcstatus <= #TCQ 0;
    end
    
  end endgenerate // end if (VC == 1)
  // }}} end VC Status Generator

  // {{{ Status Generator
  reg [CG_CTR_WIDTH-1:0]  buf_stat_codegroups_ctr;
  wire                    buf_stat_inserted;
  reg                     buf_stat_codegroups_trained_max;
  reg                     buf_stat_codegroups_lw2_max;
  reg                     buf_stat_codegroups_lw4_max;

  // The buf_stat counter expires when it reaches it 1024 codegroups this
  // varies based on the link width. Since this signal requires a a little bit
  // of time to proigate and the control symbol be generated we need to
  // provide a little leeway from 1024 to generate the signal in time.
  // If a ccomp sequence is request at the same time, we need to give enough
  // time to finish the ccomp sequence and propigate this request as well.
  // This will cost a few more cycles, so to pick a safe number of time, 15
  // cycles leeway is used.
  localparam BUF_STAT_LEEWAY      = 20;
  localparam BUF_STAT_MAX_TRAINED = 128-BUF_STAT_LEEWAY;
  localparam BUF_STAT_MAX_LW2     = 256-BUF_STAT_LEEWAY;
  // x4 needs extra time since latency is added though the OPLM due to the OPLM being a 
  // 128-bit interface only in x4 mode
  localparam BUF_STAT_MAX_LW4     = 512-BUF_STAT_LEEWAY-6;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      buf_stat_codegroups_trained_max <= #TCQ 0;
      buf_stat_codegroups_lw2_max     <= #TCQ 0;
      buf_stat_codegroups_lw4_max     <= #TCQ 0;
    end else begin
      if (!buf_stat_int_expired || buf_stat_inserted) begin
        buf_stat_codegroups_trained_max <= #TCQ (buf_stat_codegroups_ctr == BUF_STAT_MAX_TRAINED-1);
        buf_stat_codegroups_lw2_max     <= #TCQ (buf_stat_codegroups_ctr == BUF_STAT_MAX_LW2-1);
        buf_stat_codegroups_lw4_max     <= #TCQ (buf_stat_codegroups_ctr == BUF_STAT_MAX_LW4-1);
      end
    end
  end

  wire buf_stat_trained_max = PP_mode_1x && buf_stat_codegroups_trained_max;

  // For a x1 core the counter will count to 128 to meet this requirement
  // w/15 cycles of leeway, compare to 118
  generate if (LINK_WIDTH == 1) begin: buf_stat_exp_gen_x1
    assign buf_stat_int_expired = buf_stat_codegroups_trained_max;

  // For a x2 core the counter will count to 256 to meet this requirement
  // w/15 cycles of leeway, compare to 241
  end else if (LINK_WIDTH == 2) begin: buf_stat_exp_gen_x2
    assign buf_stat_int_expired = buf_stat_codegroups_lw2_max || buf_stat_trained_max;
  
  // For a x4 core the counter will count to 512 to meet this requirement
  // w/15 cycles of leeway, compare to 497. 20 is used incase a clk comp
  // request occurs when the status needs to go out.
  end else if (LINK_WIDTH == 4) begin: buf_stat_exp_gen_x4
    assign buf_stat_int_expired = buf_stat_codegroups_lw4_max || buf_stat_trained_max;
  end endgenerate

  //*COVERAGE*
  //(cp_stat_exp_w_ccomp_seq_idle1): See the buf status insertion expire at the same time a ccomp sequence 
  //is requested in idle1

  //*COVERAGE*
  //(cp_stat_exp_w_ccomp_seq_idle2): See the buf status insertion expire at the same time a ccomp sequence 
  //is requested in idle1

  //*COVERAGE*
  //(cp_buf_stat_int_expired): Cover the buf status insertion interval expires (buf_stat_int_expired).

  //*COVERAGE*
  //(cp_buf_stat_expires_before_link_init): Cover the buf status insertion
  //interval expires before the link has initialized.

  //*ASSERTION*
  //(ap_embed_buf_stat): If the buf_stat insertion interval expires, embed
  //must assert with send_status

  // A status, pa, pr functions all include the buf_status field
  assign buf_stat_inserted = (ack_status || ack_pa || ack_pr);
 
  // The Codegroups counter determines how many codegroups have been sent for
  // this link width. A VC Status must be sent every 1024-codegroups only after
  // the port initialized
  // REQ: req_pt_buf_stat_sent_every_1024
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      buf_stat_codegroups_ctr <= #TCQ 0;
    end else begin
      if (buf_stat_inserted || !PP_port_initialized) begin
        buf_stat_codegroups_ctr <= #TCQ 0;
      
      // Hold value at the max so that the status symbol will be embeded
      end else if (!buf_stat_int_expired) begin
        buf_stat_codegroups_ctr <= #TCQ buf_stat_codegroups_ctr + 1'b1;
      end
    end
  end

  //*ASSERTION*
  //(ap_buf_stat_ctr_rollover): The buffer status cg counter does not rollover

  // Send the status symbol if:
  // 1. the init_seq_ctr indicates to
  // 2. the status counter expires
  // 3. we just sent an lresp and are in tx flow control mode

  assign send_status = (send_status_init_seq || buf_stat_int_expired || lresp_sent_send_stat) && 
                       !buf_stat_inserted;
  // }}} end Status Generator
 
  // {{{ Stype1 Function Generator
  // The stype1 generator generates stype1 functions with the 
  // following priority:
  // 1. LREQ-reset-device from UG  
  // 2. LREQ-input-status from OLLM RX
  // 3. MCE (multicast-event)
  // 4. RFR (restart-from-retry)
  // 5. SOP (start-of-packet)
  // 6. EOP (end-of-packet)
  // 7. LREQ-any from PHY CFG 
  // 8. NOP (always the default)
  
  // When a LREQ arrives from the config latch the request since it is only one
  // cycle
  reg       lreq_cfg;
  reg [2:0] lreq_cmd_cfg;
  wire      send_lreq_cfg;

  // Mask off the lreq if there is already one outstanding
  assign in_packet = PTA_in_packet || PTB_in_packet;

  assign send_lreq_cfg = lreq_cfg && !PR_output_error_stop && !ack_lreq && 
                         !in_packet;
  
  //Ask a LREQ request from the phy config whenever one is sent with the same
  //command.  This way if the two requests with the same command occur, only one will
  //be sent.
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      lreq_cfg     <= #TCQ 0;
      lreq_cmd_cfg <= #TCQ 0;
    end else begin
      // Mask off all LREQs from the config space if the port is not
      // initialized.
      if (PC_send_lreq && PP_port_initialized) begin
        lreq_cfg     <= #TCQ 1'b1;
        lreq_cmd_cfg <= #TCQ PC_lreq_cmd;

      end else if (ack_lreq) begin
        lreq_cfg     <= #TCQ 0;
        lreq_cmd_cfg <= #TCQ 0;
      end
    end
  end

  // When an MCE arrives from the user latch it in case it needs to be stalled
  // for link_initialization
  reg mce_request;

  //Ack an MCE when it has been inserted
  assign ack_mce = (stype1_0_mce || stype1_1_mce) && PTR_pts_advance;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PTS_mce_sent <= #TCQ 0;
    end else begin
      PTS_mce_sent <= #TCQ ack_mce;
    end
  end

  //Send the MCE only if the link is initialized
  wire send_mce = mce_request && !ack_mce;
  wire send_stomp_1 = PTB_src_disc; // cr 800810, stomp

  reg send_stomp_d;
  wire send_stomp;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      send_stomp_d <= #TCQ 1'b0;
    end else begin
      send_stomp_d <= #TCQ send_stomp_1;
    end
  end
  assign send_stomp = send_stomp_d || send_stomp_1;// cr 800810, stomp

  // CROSS Clock domain here. This is intentionally asynchronous.
  reg [1:0] ug_phy_mce_srl;
  reg       ug_phy_mce_q, ug_phy_mce_qq;
  always @(posedge phy_clk or posedge UG_phy_mce) begin
    if (UG_phy_mce) begin
      ug_phy_mce_srl <= #TCQ 2'b11;
    end else if (phy_rst_q) begin
      ug_phy_mce_srl <= #TCQ 2'b00;
    end else begin
      ug_phy_mce_srl <= #TCQ {ug_phy_mce_srl[0], 1'b0};
    end
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      ug_phy_mce_q  <= #TCQ 1'b0;
      ug_phy_mce_qq <= #TCQ 1'b0;
    end else begin
      ug_phy_mce_q  <= #TCQ |ug_phy_mce_srl;
      ug_phy_mce_qq <= #TCQ ug_phy_mce_q;
    end
  end


  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      mce_request <= #TCQ 0;
    end else begin
      // Check to see that a new MCE is not asserted on the same cycle one
      // was sent, if so dont drop mce_request until another is sent.
      if (ack_mce && !(ug_phy_mce_q && !ug_phy_mce_qq)) begin
        mce_request <= #TCQ 0;

      end else if (ug_phy_mce_q && !ug_phy_mce_qq && PR_link_initialized) begin
        mce_request <= #TCQ 1;
      end
    end
  end

  // Send a link reset as long as PTB_link_reset is asserted
  // Register it in case it is only asserted for one cycle, one will still be
  // sent.
  wire ack_lreq_rd = (stype1_0_lreq_rd) && PTR_pts_advance;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      link_reset_request <= #TCQ 0;
    end else begin
      // Check to see that a new MCE is not asserted on the same cycle one
      // was sent, if so dont drop mce_request until another is sent.
      if (!PTB_link_reset) begin
        link_reset_request <= #TCQ 0;

      end else if (!PR_send_lreq) begin
        link_reset_request <= #TCQ 1;
      end
    end
  end

  always @* begin
    send_link_reset = link_reset_request && !in_packet;
  end

  //*COVERAGE*
  //(cp_lreq_reset_w_ollmrx_is): See a link reset occur when the ollm rx requests an 
  // input status to be sent
 
  //*COVERAGE*
  //(cp_link_reset_w_ccomp): See a link reset collisions with a ccomp request
  
  // Sort the stype1 function according to there priority left to right
  
  // Overwrite the eop with an sop if another packet is being sent b2b to the
  // current packet and there does not need to be a break inserted for the
  // ccomp_sequence
  // REQ: req_pt_completed_pkt_ended_correctly
  // REQ: req_pt_killed_pkt_ended_correctly
  reg  send_overwrite_sop;
  reg  send_overwrite_sop_q;
  reg  send_starting_sop;
  reg  send_starting_sop_q;
  wire kill_queued_eop;
  reg  send_ending_eop;

  wire ack_sop = stype1_sop && PTR_pts_advance;

  wire single_cycle = PTB_sop && PTB_eop;
  
  // Do not override an EOP if we need to send the ccomp sequence.
  // Override the EOP with an SOP if we see an SOP coming. This can occur from
  // the assertion of PTB_sop_d, except if in the case of a clk comp we need
  // to look at PTB_sop since we know the data mux is stalling PTA on an
  // SOP already.
  wire overwrite_sop = (PTB_sop_d && PTB_eop && PTR_ptb_advance);

  // Queue up SOP requests when:
  // 1. We are at the start of a packet
  // 2. We are in need of both an overwrite SOP plus another SOP in the case
  //    of a single cycle packet
  // For overrides only advance if pta advance is asserted so the cs is ready
  // on eop
  // For starting sop's only advance if the buf module is advanceing
  // Timing for this is such that it lines up for the data mux 
  wire starting_sop = (PTB_sop && !send_overwrite_sop_q && PTR_pta_advance) ||
                      (single_cycle && PTB_sop_d && PTR_ptb_advance && 
                       !PP_idle2_selected && !ack_sop);

  // Clear any queued SOPs if:
  // 1. A starting SOP is acked
  always @* begin
    if (ack_sop && send_starting_sop_q && !(overwrite_sop && send_overwrite_sop_q)) begin 
      send_starting_sop = 1'b0;
    end else if (starting_sop) begin
      send_starting_sop = 1'b1;
    end else begin
      send_starting_sop = send_starting_sop_q;
    end
  end

  // Queue up SOP requests for when we are overwritting an EOP
  // Kill an override if: 
  // 1. Kill an overriding SOP for a non-single cycle pkt when the last EOP is
  //    seen
  // 2. Because a single cycle pkt causes both starting_sop and overwrite sop
  //    to trigger. we need to kill the overriding sop only when the last eop is
  //    seen and the starting sop was already inserted in order to align control
  //    symbols correctly.
  wire kill_queued_sop = (send_overwrite_sop_q && PTB_eop && !PTB_sop_d && 
                          !PTB_sop && PTR_ptb_advance);
  
  always @* begin
    if (kill_queued_sop) begin
      send_overwrite_sop = 1'b0;
    end else if (overwrite_sop) begin
      send_overwrite_sop = 1'b1;
    end else if (ack_sop && send_overwrite_sop_q && !send_starting_sop_q) begin
      send_overwrite_sop = 1'b0;
    end else begin
      send_overwrite_sop = send_overwrite_sop_q;
    end
  end

  // Latch the send SOP signals
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      send_starting_sop_q  <= #TCQ 0;
      send_overwrite_sop_q <= #TCQ 0;
    end else begin
      send_starting_sop_q  <= #TCQ send_starting_sop;
      send_overwrite_sop_q <= #TCQ send_overwrite_sop;
    end
  end

  // Assert to send an SOP for either a SOP or overwriting EOP with an SOP condition
  always @* begin
    send_sop = (send_starting_sop || send_overwrite_sop) && !send_ccomp_eop;
  end

  // *COVERAGE*
  // (cr_ccomp_req_w_sop): Cover the clk compensation is request on
  // a start of packet for both a starting sop and overwriting sop
  
  //*COVERAGE*
  //(cp_link_reset_w_ccomp): See a link reset end collisions with a ccomp request
  
  //Only send an eop if we are not sending an sop on the same cycle
  //Or if there was a single cycle pkt that is ending

  reg send_ending_eop_q;
  reg single_cycle_q;

  assign ack_eop = stype1_eop && PTR_pts_advance;

  assign ending_eop = PTB_eop && PTR_ptb_advance;

  // If an EOP is killed register it so we know is an actually EOP is then 
  // needed after the killed one.
  reg queue_eop;

  // Kill a pending EOP if:
  // 1. an SOP comes with enough time to make it b2b. This will occur if the SOP arrives
  // late after an EOP is seen with no starting packet to follow.
  assign kill_queued_eop = PTS_eop && !PTR_pts_advance && send_sop && !PP_ccomp_req;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      queue_eop <= #TCQ 0;
    end else begin
      queue_eop <= #TCQ (kill_queued_eop && ending_eop && !PTB_sop_d); 
    end
  end
  

  always @* begin
    if ((queue_eop || ending_eop) && (!send_overwrite_sop || !PTB_sop_d)) begin
      send_ending_eop = 1'b1;
    end else if (ack_eop && !single_cycle_q) begin
      send_ending_eop = 1'b0;
    end else begin
      send_ending_eop = send_ending_eop_q;
    end
  end

  // latch the send_eop signal
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      send_ending_eop_q <= #TCQ 0;
    end else begin
      send_ending_eop_q <= #TCQ send_ending_eop;
    end
  end

  //latch the single_cycle signal
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      single_cycle_q <= #TCQ 0;
    end else begin
      single_cycle_q <= #TCQ single_cycle && PTR_ptb_advance;
    end
  end

  // When a ccomp_eop is pending and a new eop arrives we need to save this to
  // be sent following the ack of the ccomp_eop
  reg pending_eop_during_ccomp;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      pending_eop_during_ccomp <= #TCQ 0;
    end else begin
      if (ack_eop && !send_ccomp_eop_q) begin
        pending_eop_during_ccomp <= #TCQ 0;
      end else if (ending_eop && send_ccomp_eop_q && !PTB_sop_d) begin
        pending_eop_during_ccomp <= #TCQ 1;
      end
    end
  end

  // Indicate to send an EOP only when there is one queued up and 
  // we are not sending an SOP
  always @* begin
    send_eop = (send_ending_eop || (pending_eop_during_ccomp && !ack_eop)) && 
               !send_sop && !send_ccomp_eop;
  end

  // Figure out when to send a EOP because the ccomp sequence needing a break
  // in the transmit stream
  reg pta_in_packet_q;

  // Do not grant the ccomp sequence until any pending MCEs are sent to get
  // them out quickly.
  always @* begin
    if (ack_eop) begin
      send_ccomp_eop = 0;
    end else if (PP_ccomp_req && ending_eop && pta_in_packet_q && PTA_in_packet && !mce_request) begin
      send_ccomp_eop = 1;
    end else begin
      send_ccomp_eop = send_ccomp_eop_q;
    end
  end

  //latch the send ccomp_eop and pta_in_packet signals
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      send_ccomp_eop_q <= #TCQ 0;
      pta_in_packet_q  <= #TCQ 0;
    end else begin
      send_ccomp_eop_q <= #TCQ send_ccomp_eop;
      pta_in_packet_q  <= #TCQ PTA_in_packet;
    end
  end
  
  //*ASSERTION*
  //(ap_sop_and_eop_generated): sop and eop cannot occur on the same cycle for
  //IDLE1 mode.

  //REQ: req_pt_stype1_cs_priorities
  //REQ: req_pt_mce_minimal_latency
  
  //Only queue up a cs if it wasnt just sent
  assign send_lreq = (PR_send_lreq && !PTS_lreq_sent) && !ack_lreq && !in_packet;
  assign send_rfr  = (PR_send_rfr && !PTS_rfr_sent) && !ack_rfr && !in_packet;

  wire [7:0] stype1_functions_0 = {send_mce, send_ccomp_eop, send_sop, send_eop, 
                                   send_link_reset, send_rfr, send_lreq, send_lreq_cfg};

  //*COVERAGE* 
  //(cr_stype1_functions_0): Cross PTB_link_reset, send_mce, with PTA_in_packet
 
  //*COVERAGE*
  //(cp_lreq): An lreq occurs from the PHY config and the OLLM RX as well as
  //independently

  //*COVERAGE*
  //(cp_two_reset_device_lreqs_occur): PTB_link_reset and send_lreq_cfg
  //with lreq_cmd_cfg == RESET_DEVICE_CMD occurs.

  //*COVERAGE*
  //(cp_two_input_status_lreqs_occur): PR_send_lreq and send_lreq_cfg
  //with lreq_cmd_cfg == INPUT_STATUS_CMD occurs.
 
  //*COVERAGE*
  //(cp_resetdevice_user_w_inputstatus_cfg): See a reset device from the user with a
  //input status request from the config at the same time

  //*COVERAGE*
  //(cp_rfr_killed_pkt_on_eop, cp_lreq_killed_pkt_on_eop, 
  // cp_lreq_killed_pkt_mid_pkt, cp_rfr_killed_pkt_mid_pkt):
  // Cover a packet is killed with a RFR and an LREQ with and without EOP being asserted.

  //*COVERAGE*
  //(cp_overwrite_eop_w_ccompreq): Cover an overwrite condition needs to take
  //place at the same time a clk compensation sequence is requested.

  //*COVERAGE*
  //(cp_ccompreq_X_sop): Cross ccomp_req with an SOP

  //*COVERAGE*
  //(cp_ccompreq_X_eop): Cross ccomp_req with an EOP
  
  // Get the one hot version of the function to send
  assign stype1_onehot_0 = stype1_onehot(stype1_functions_0);
  // Get the binary version of the function 
  assign stype1_binary_0 = stype1_binary(stype1_functions_0);

  // Only generate a new symbol if:
  // 1. No symbol is currently valid and there isnt one that is trying to be
  //    embedded from an stype0 unless its the end of a packet already. This
  //    is because it may try to embed a packet delimiting control symbol
  //    incorrectly otherwise.
  // 2. The valid one has been accepted
  // 4. An SOP is killed and needs to be replaced with an EOP
  wire advance_stype1 = (!stype1_valid_0 && (!stype0_embed_0 || (PTA_eop && PTR_pta_advance))) || 
                         PTR_pts_advance || kill_queued_sop || kill_queued_eop;
  // Generate the embed flag with the symbol
  // Need to force the symbol if 
  // 1. we are sending a multicast event control symbol
  // REQ: req_pt_no_invalid_cs_in_pkt
  wire stype1_embed_req_0 = stype1_onehot_0[MCE_BIT];

  // Based on the selected stype1, generate the function fields
  // REQ: req_pt_cs_pd_delimiter_used_correctly
  // REQ: req_pt_cs_sc_delimiter_used_correctly
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      delimiter_0      <= #TCQ SC;
      stype1_cmd_0     <= #TCQ NO_CMD;
      stype1_0         <= #TCQ STYPE1_NOP;
      stype1_valid_0   <= #TCQ 0;
      stype1_embed_0   <= #TCQ 0;
      stype1_0_mce     <= #TCQ 0;
      stype1_0_rfr     <= #TCQ 0;
      stype1_0_lreq    <= #TCQ 0;
      stype1_0_lreq_rd <= #TCQ 0;
    end else begin
      if (advance_stype1) begin
        delimiter_0      <= #TCQ stype1_delimiter(stype1_binary_0);
        stype1_cmd_0     <= #TCQ stype1_cmd(stype1_binary_0,lreq_cmd_cfg);
        stype1_0         <= #TCQ stype1_type(stype1_binary_0);
	  //enable below line and comment above line for stype_1_0 logic in case the STOMP functionality is decided to be added 
      //stype1_0         <= #TCQ send_stomp? 3'b001:stype1_type(stype1_binary_0);//  cr 800810, stomp
	    //stype1_0         <= #TCQ send_stomp_1? 3'b001:stype1_type(stype1_binary_0);// dont un comment this line
        stype1_valid_0   <= #TCQ |stype1_onehot_0; 
        stype1_embed_0   <= #TCQ stype1_embed_req_0;

        // Save off the type of control symbol to improve timing 
        stype1_0_mce     <= #TCQ stype1_onehot_0[MCE_BIT];
        stype1_0_rfr     <= #TCQ stype1_onehot_0[RFR_BIT];
        stype1_0_lreq    <= #TCQ stype1_onehot_0[LREQ_USERDEF_BIT] ||
                                 stype1_onehot_0[LREQ_INPUT_STATUS_BIT];
        stype1_0_lreq_rd <= #TCQ stype1_onehot_0[LREQ_RESET_DEVICE_BIT];                     
      end
    end
  end

  // Only generate a second stype1 function if IDLE1 mode is possible
  generate if (IDLE1) begin: stype1_1_gen
    reg [7:0] stype1_functions_1;

    always @* begin
      // Since we need LREQ/reset-device's to be back to back exiting the core
      // IDLE1 is special in that it needs to generate two per cycle to fill
      // the 4 byte GT interface. So this special case handles generating
      // a LREQ/reset only when stype _0 is a LREQ/reset
      if (stype1_onehot_0[LREQ_RESET_DEVICE_BIT]) begin
        // mask the LREQ/reset if another stype is going out
        stype1_functions_1 = LREQ_RESET_DEVICE_ONEHOT;

      // Get the new one hot for the second symbol omiting the the symbol on the
      // *_0 fields and masking sending a reset device unless it has started
      // being sent
      end else begin
        stype1_functions_1 = (stype1_functions_0 ^ stype1_onehot_0) & 8'b1111_1011;
      end
    end
    
    // Get the onehot/binary encoding for the stype1 second function
    assign stype1_onehot_1 = stype1_onehot(stype1_functions_1);
    assign stype1_binary_1 = stype1_binary(stype1_functions_1);

    // Generate the embed flag with the symbol
    // Need to force the symbol if 
    // 1. we are sending a multicast event control symbol
    // REQ: req_pt_no_invalid_cs_in_pkt
    wire stype1_embed_req_1 = stype1_onehot_1[MCE_BIT];
    
    // Based on the selected stype1, generate the function fields for the 
    // second control symbol
    always @(posedge phy_clk) begin
      if (phy_rst_q) begin
        delimiter_1     <= #TCQ SC;
        stype1_cmd_1    <= #TCQ NO_CMD;
        stype1_1        <= #TCQ STYPE1_NOP;
        stype1_valid_1  <= #TCQ 0;
        stype1_embed_1  <= #TCQ 0;
        stype1_1_mce    <= #TCQ 0;
        stype1_1_rfr    <= #TCQ 0;
        stype1_1_lreq   <= #TCQ 0;
        
      // Only generate a second control symbol if not in IDLE2 mode
      end else if (!PP_idle2_selected) begin
        if (advance_stype1) begin
          delimiter_1     <= #TCQ stype1_delimiter(stype1_binary_1);
          stype1_cmd_1    <= #TCQ stype1_cmd(stype1_binary_1,lreq_cmd_cfg);
          stype1_1        <= #TCQ stype1_type(stype1_binary_1);
          stype1_valid_1  <= #TCQ |stype1_onehot_1;
          stype1_embed_1  <= #TCQ stype1_embed_req_1;

          // Save off the type of control symbol to improve timing
          stype1_1_mce    <= #TCQ stype1_onehot_1[MCE_BIT];
          stype1_1_rfr    <= #TCQ stype1_onehot_1[RFR_BIT];
          stype1_1_lreq   <= #TCQ stype1_onehot_1[LREQ_USERDEF_BIT] ||
                                  stype1_onehot_1[LREQ_INPUT_STATUS_BIT] ||
                                  stype1_onehot_1[LREQ_RESET_DEVICE_BIT];
        end
      end
    end

  //*ASSERTION*
  //(ap_rogue_stype1_embed_0): stype1_embed_0 can not assert with no valid control symbols

  //*ASSERTION*
  //(ap_rogue_stype1_embed_1): stype1_embed_1 can not assert with no valid control symbols

  // Tie off the onehot_1 signal when IDLE1 is not set
  end else begin: no_stype1_1_gen
    always @(posedge phy_clk) begin
      stype1_cmd_1  <= #TCQ NO_CMD;
      stype1_1      <= #TCQ STYPE1_NOP;
      stype1_1_rfr  <= #TCQ 0;
      stype1_1_lreq <= #TCQ 0;
      stype1_1_mce  <= #TCQ 0;
    end

    assign stype1_onehot_1 = 0;
    assign stype1_binary_1 = 0;
  end endgenerate //end if (IDLE1)

  // Create a register SOP and EOP signal to improve timing
  generate 
    case ({(IDLE1 == 1),(IDLE2 == 1)})
      //IDLE1 Only
      {1'b1,1'b0}: begin: idle1_sop_eop_gen
        always @(posedge phy_clk) begin
          if (phy_rst_q) begin
            stype1_sop <= #TCQ 0;
            stype1_eop <= #TCQ 0;
          end else begin
            if (advance_stype1) begin
              stype1_sop <= #TCQ stype1_onehot_0[SOP_BIT] || stype1_onehot_1[SOP_BIT];
              stype1_eop <= #TCQ stype1_onehot_0[EOP_BIT] || stype1_onehot_0[CCOMP_EOP_BIT] ||
                                 stype1_onehot_1[EOP_BIT] || stype1_onehot_1[CCOMP_EOP_BIT];
            end
          end 
        end
      end 

      // IDLE2 Only
      {1'b0,1'b1}: begin: idle2_sop_eop_gen
        always @(posedge phy_clk) begin
          if (phy_rst_q) begin
            stype1_sop <= #TCQ 0;
            stype1_eop <= #TCQ 0;
          end else begin
            if (advance_stype1) begin
              stype1_sop <= #TCQ stype1_onehot_0[SOP_BIT];
              stype1_eop <= #TCQ stype1_onehot_0[EOP_BIT] || stype1_onehot_0[CCOMP_EOP_BIT];
            end
          end 
        end
      end

      // IDLE1 and IDLE2
      {1'b1,1'b1}: begin: idle2_sop_eop_gen
        always @(posedge phy_clk) begin
          if (phy_rst_q) begin
            stype1_sop <= #TCQ 0;
            stype1_eop <= #TCQ 0;
          end else begin
            if (advance_stype1) begin
              stype1_sop <= #TCQ (PP_idle2_selected) ? 
                                  stype1_onehot_0[SOP_BIT] :
                                  (stype1_onehot_0[SOP_BIT] || stype1_onehot_1[SOP_BIT]);
              stype1_eop <= #TCQ (PP_idle2_selected) ?
                                  (stype1_onehot_0[EOP_BIT] || stype1_onehot_0[CCOMP_EOP_BIT]) :
                                  (stype1_onehot_0[EOP_BIT] || stype1_onehot_0[CCOMP_EOP_BIT] ||
                                   stype1_onehot_1[EOP_BIT] || stype1_onehot_1[CCOMP_EOP_BIT]);
            end
          end 
        end
      end //end idle2 only
    endcase
  endgenerate //end sop/eop generation

  //*ASSERTION*
  //(ap_invalid_stype1_valid): Valid can not be asserted on stype1_valid_1
  //without a valid on stype1_valid_0

  // Acknowledge control symbol requests if they were requested by the OLLM RX
  assign ack_lreq = (stype1_0_lreq || stype1_1_lreq) && PTR_pts_advance;
  assign ack_rfr  = (stype1_0_rfr || stype1_1_rfr) && PTR_pts_advance;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PTS_lreq_sent   <= #TCQ 0;
      PTS_rfr_sent    <= #TCQ 0;
    end else begin
      PTS_lreq_sent   <= #TCQ ack_lreq && PR_send_lreq;
      PTS_rfr_sent    <= #TCQ ack_rfr && PR_send_rfr;
    end
  end 

  // {{{ + STYPE1 Utility Functions +
  // {{{ stype1_delimiter -
  // returns the delimiter for the stype1 function
  wire eop_accepted = PTS_eop && PTR_pts_advance;

  function [7:0] stype1_delimiter (
    input [3:0] functions
  ); begin
      case (functions)
        SOP_BINARY,EOP_BINARY, CCOMP_EOP_BINARY: stype1_delimiter = PD;
        default:                                 stype1_delimiter = SC;
      endcase
    end 
  endfunction
  // }}} end stype0_cmd

  // {{{ stype1_cmd -
  // returns the cmd feild for the stype1 function
  function [2:0] stype1_cmd (
    input [3:0] functions,
    input [2:0] lreq_cmd_cfg
  ); begin
      case (functions)
        LREQ_RESET_DEVICE_BINARY:     stype1_cmd = RESET_DEVICE_CMD;
        LREQ_INPUT_STATUS_BINARY:     stype1_cmd = INPUT_STATUS_CMD;
        LREQ_USERDEF_BINARY:          stype1_cmd = lreq_cmd_cfg;
        default:                      stype1_cmd = NO_CMD;
      endcase
    end 
  endfunction
  // }}} end stype0_cmd
  
  // {{{ stype1_type -
  // returns the stype1 type feild for an stype1 function
  function [2:0] stype1_type (
    input [3:0] functions
  ); begin
      case (functions)
        LREQ_RESET_DEVICE_BINARY:     stype1_type = STYPE1_LREQ;
        LREQ_INPUT_STATUS_BINARY:     stype1_type = STYPE1_LREQ;
        MCE_BINARY:                   stype1_type = STYPE1_MCE;
        RFR_BINARY:                   stype1_type = STYPE1_RFR;
        SOP_BINARY:                   stype1_type = STYPE1_SOP;
        EOP_BINARY, CCOMP_EOP_BINARY: stype1_type = STYPE1_EOP;
        LREQ_USERDEF_BINARY:          stype1_type = STYPE1_LREQ;
        NOP_BINARY:                   stype1_type = STYPE1_NOP;
        default:                      stype1_type = {3{1'bX}};
      endcase
    end 
  endfunction
  // }}} end stype1_type

  // {{{ stype1_onehot -
  // returns the one hot encoding of the valid stype1 functions
  function [7:0] stype1_onehot (
    input [7:0] functions
  ); begin
      casex ({functions})
        {8'b1xxx_xxxx}: stype1_onehot = MCE_ONEHOT;        
        {8'b01xx_xxxx}: stype1_onehot = CCOMP_EOP_ONEHOT;        
        {8'b001x_xxxx}: stype1_onehot = SOP_ONEHOT;
        {8'b0001_xxxx}: stype1_onehot = EOP_ONEHOT;
        {8'b0000_1xxx}: stype1_onehot = LREQ_RESET_DEVICE_ONEHOT;
        {8'b0000_01xx}: stype1_onehot = RFR_ONEHOT;
        {8'b0000_001x}: stype1_onehot = LREQ_INPUT_STATUS_ONEHOT;
        {8'b0000_0001}: stype1_onehot = LREQ_USERDEF_ONEHOT;
        {8'b0000_0000}: stype1_onehot = NOP_ONEHOT;
        default       : stype1_onehot = {7{1'bX}};
      endcase
    end 
  endfunction
  // }}} end stype1_onehot

  // {{{ stype1_binary -
  // returns the binary encoding of the valid stype1 functions
  function [3:0] stype1_binary (
    input [7:0] functions
  ); begin
      casex ({functions})
        {8'b1xxx_xxxx}: stype1_binary = MCE_BINARY;        
        {8'b01xx_xxxx}: stype1_binary = CCOMP_EOP_BINARY;        
        {8'b001x_xxxx}: stype1_binary = SOP_BINARY;
        {8'b0001_xxxx}: stype1_binary = EOP_BINARY;
        {8'b0000_1xxx}: stype1_binary = LREQ_RESET_DEVICE_BINARY;
        {8'b0000_01xx}: stype1_binary = RFR_BINARY;
        {8'b0000_001x}: stype1_binary = LREQ_INPUT_STATUS_BINARY;
        {8'b0000_0001}: stype1_binary = LREQ_USERDEF_BINARY;
        {8'b0000_0000}: stype1_binary = NOP_BINARY;
        default       : stype1_binary = {4{1'bX}};
      endcase
    end 
  endfunction
  // }}} end stype1_binary

  // }}} + STYPE0 Utility Functions +
  // }}} end Stype1 Function Generator

  // {{{ + Short Control Symbol Creation +
  // Only generate support for short control symbols if IDLE1 is set
  //REQ: req_pt_short_cs_idle1
  //REQ: req_pt_no_short_cs_idle1_disabled
  generate if (IDLE1) begin: short_cs_gen
    // Concatinate the fields together to form the cs fields for a short
    // control symbol
    // Only grab 5-bits of the parameter fields in case that IDLE2 is set
    // and the default widths are 6-bits the parameters
    // REQ: req_pt_cs_functions_are_packed
    wire [18:0] short_cs_fields_0 = {stype0_0, parameter0_0[4:0], parameter1_0[4:0], 
                                     stype1_0, stype1_cmd_0};
    wire [18:0] short_cs_fields_1 = {stype0_1, parameter0_1[4:0], parameter1_1[4:0], 
                                     stype1_1, stype1_cmd_1};

    //*COVERAGE*
    //(cr_all_stypes): cover all combinations of stype0_0, stype0_1,
    //stype1_0, stype1_1

    //*ASSERTION*
    //(ap_idle1_cs_param0_invalid): For both IDLE1 and IDLE2 mode, if PP_idle2_selected is low 
    //the parameter fields bit[5] must be 0.

    //*ASSERTION*
    //(ap_idle1_cs_param1_invalid): For both IDLE1 and IDLE2 mode, if PP_idle2_selected is low 
    //the parameter fields bit[5] must be 0.
  
    // Use the cs fields to generate the 5-bit CRC
    wire [4:0] cs_fields_0_crc5;
    wire [4:0] cs_fields_1_crc5;
 
    //REQ: req_pt_crc5_correct_bits_used
    srio_gen2_v4_1_16_crc5_20 short_crc_cs0_inst (
      .crc    (cs_fields_0_crc5),
      .din    (short_cs_fields_0));

    srio_gen2_v4_1_16_crc5_20 short_crc_cs1_inst (
      .crc    (cs_fields_1_crc5),
      .din    (short_cs_fields_1));
    
    //REQ: rreq_pt_cs_delimited
    //REQ: req_pt_short_cs_delimited
    //REQ: req_pt_short_cs_crc5
    wire [31:0] control_symbol_0 = {delimiter_0, short_cs_fields_0, cs_fields_0_crc5};
    wire [31:0] control_symbol_1 = {delimiter_1, short_cs_fields_1, cs_fields_1_crc5};

    // Add the delimiter and CRC
    assign short_cs_data  = {control_symbol_0, control_symbol_1};
    assign short_cs_valid = {(stype0_valid_0 | stype1_valid_0), stype1_valid_1};
    assign short_cs_embed = stype0_embed_0 | stype1_embed_0 | stype1_embed_1;

    // Only the delimiters are K characters this can be tied off since it will
    // be masked with valid
    assign short_cs_charisk  = 8'b1000_1000;

    // Do not use the lreq field for IDLE1 mode
    assign short_cs_lreq  = 0;

    assign short_cs_sop = stype1_sop;
    assign short_cs_eop = stype1_eop;

    //*COVERAGE*
    //(cr_stype0_X_stype1): cross stype0_valid_0, stype1_valid_0, stype1_valid_1
    //It is not legal for {stype1_valid_0, stype1_valid_1} == 2'b01

    //*ASSERTION*
    //(ap_short_embedded): If short_cs_embed is asserted, stype1_0 and stype1_1
    //must be a MCE or NOP
    
    // Stall if two control symbols are generated and a full dword of packet
    // data is coming, this will cause the packet data to stall an extra cycle
    // first so the two cs's can be inseterted. This only needs to occur when 
    // we are out of packet because the data mux will handle the case when we
    // are in packet.
    wire two_cs = (|stype1_binary_0 && |stype1_binary_1); 

    wire sop_next = (stype1_onehot_0[SOP_BIT] || stype1_onehot_1[SOP_BIT]);

    always @(posedge phy_clk) begin
      if (phy_rst_q) begin
        short_cs_stall <= #TCQ 0;
      end else begin
        if (PTR_pts_advance || !(&PTA_valid_d)) begin
          short_cs_stall <= #TCQ two_cs && &PTA_valid_d && PTR_ptb_advance && 
                                 (!PTA_in_packet || (PTA_in_packet && PTR_pts_advance && sop_next));
      
        end
      end
    end

  end endgenerate //if (IDLE1)
  // }}} + end Short Control Symbol Creation +
  
  // {{{ + Long Control Symbol Creation +
  // REQ: req_pt_no_long_cs_idle2_disabled
  generate if (IDLE2) begin: long_cs_gen
    // Concatinate the fields together to form the cs fields for a long control
    // symbol
    // Only use the fields from *_0 since it will take the entire 64-bit bus.
    // REQ: req_pt_cs_functions_are_packed
    wire [34:0] long_cs_fields = {stype0_0, parameter0_0, parameter1_0, 
                                  stype1_0, stype1_cmd_0, 14'b0};

    // Use the cs fields to generate the 13-bit CRC
    wire [12:0] cs_fields_crc13;
    
    srio_gen2_v4_1_16_crc13_35 long_cs_inst (
      .crc    (cs_fields_crc13),
      .din    (long_cs_fields));  
    
    // Add the delimiter and CRC
    //REQ: req_pt_long_cs_idle2
    //REQ: rreq_pt_cs_delimited
    //REQ: req_pt_long_cs_start_delimiter
    //REQ: req_pt_long_cs_end_delimiter
    //REQ: req_pt_long_cs_start_eq_end_delimiter
    assign long_cs_data  = {delimiter_0, long_cs_fields, cs_fields_crc13, delimiter_0};
    assign long_cs_valid = {2{(stype0_valid_0 | stype1_valid_0)}};
    assign long_cs_embed = (stype0_embed_0) | (stype1_embed_0);
    assign long_cs_lreq  = (stype1_0 == STYPE1_LREQ);

    // Only the delimiters are K characters this can be tied off since it will
    // be masked with valid
    assign long_cs_charisk  = 8'b1000_0001;

    assign long_cs_sop = stype1_sop;
    assign long_cs_eop = stype1_eop;
    
    //*ASSERTION*
    //(ap_long_embedded): If long_cs_embed is asserted, stype1_0
    //must be a MCE or NOP

    // Stall data for control symbols since they will take a whole cycle to send
    always @(posedge phy_clk) begin
      if (phy_rst_q) begin
        long_cs_stall <= #TCQ 0;
      end else begin
        long_cs_stall <= #TCQ (|stype0_onehot_0 || |stype1_onehot_0) && 
                              (&PTA_valid_d && !PTA_in_packet && PTR_ptb_advance);
      end
    end

  end endgenerate //if (IDLE2)
  // }}} + end Long Control Symbol Creation +
  
  // {{{ Control Symbol Selector
  // Select the appropriate length control symbol based on the parameters
  // or the PP_idle2_selected signal
  generate case ({(IDLE2 == 1), (IDLE1 == 1)})
    // IDLE2 Only mode
    {1'b1,1'b0}: begin: idle2_only_cs_select_gen
      assign PTS_data     = long_cs_data;
      assign PTS_valid    = long_cs_valid;
      assign PTS_embed_cs = long_cs_embed;
      assign PTS_lreq     = long_cs_lreq;
      assign PTS_charisk  = long_cs_charisk;
      assign PTS_sop      = stype1_sop;
      assign PTS_eop      = stype1_eop;
      assign PTS_stall    = long_cs_stall;

    end
    // IDLE1 Only mode
    {1'b0,1'b1}: begin: idle1_only_cs_select_gen
      assign PTS_data     = short_cs_data;
      assign PTS_valid    = short_cs_valid;
      assign PTS_embed_cs = short_cs_embed; 
      assign PTS_lreq     = short_cs_lreq;
      assign PTS_charisk  = short_cs_charisk;
      assign PTS_sop      = stype1_sop;
      assign PTS_eop      = stype1_eop;
      assign PTS_stall    = short_cs_stall;
    end

    // IDLE1 and IDLE 2 modes
    {1'b1,1'b1}: begin: idle12_cs_select_gen
      assign PTS_data     = (PP_idle2_selected) ? long_cs_data    : short_cs_data;
      assign PTS_valid    = (PP_idle2_selected) ? long_cs_valid   : short_cs_valid;
      assign PTS_embed_cs = (PP_idle2_selected) ? long_cs_embed   : short_cs_embed;  
      assign PTS_lreq     = (PP_idle2_selected) ? long_cs_lreq    : short_cs_lreq;  
      assign PTS_charisk  = (PP_idle2_selected) ? long_cs_charisk : short_cs_charisk;  
      assign PTS_sop      = stype1_sop;  
      assign PTS_eop      = stype1_eop;
      assign PTS_stall    = (PP_idle2_selected) ? long_cs_stall   : short_cs_stall;
    end
  endcase endgenerate
  
  //*ASSERTION*
  //(ap_cs_lreq): cs_lreq can not assert without valid data indicated by PTS_valid

  //*ASSERTION*
  //(ap_cs_embed): cs_embed can not assert without valid data indicated by PTS_valid
  // }}} IDLE Sequence Selector  

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2010 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/phy/ollm_tx/srio_gen2_v4_1_16_ollm_tx_pkt_assembly.v#1 $
//----------------------------------------------------------------------
//
// OLLM_TX_PKT_ASSEMBLY
// Description:
// This module is responsible for accepting the packets from the 
// ollm_tx_buf_axi module and adding the ackID, CRC, and Pad
//
// Hierarchy:
// PHY_TOP
//    |___OLLM_TX_TOP
//             |_____OLLM_TX_READY_GEN
//             |_____OLLM_TX_BUF
//             |_____OLLM_TX_PKT_ASSEMBLY <-- this module
//             |_____OLLM_TX_CS_GEN
//             |_____OLLM_TX_DATA_MUX
//             |_____OLLM_TX_OPLM
// ---------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_ollm_tx_pkt_assembly
  #(
    parameter TCQ         = 100,
    parameter IDLE2       = 0,   // Include the IDLE2 Sequence {0,1}
    parameter SWITCH_MODE = 0    // Core generated with switch mode support
  )      
  (
    // {{{ Port Declarations
    // System Signals
    input               phy_clk,                // PHY interface clock
    input               phy_rst,                // Reset for PHY clock Domain
   
    // OLLM RX Interface
    output reg          PT_switch_crc_err,      // There was an error on the Final CRC

    // OLLM TX Buf AXI Interface
    input               PTB_sop,                // SOP
    input               PTB_eop,                // EOP
    input        [63:0] PTB_data,               // Data
    input        [3:0]  PTB_keep,               // Strobe
    input               PTB_valid,              // Valid Data
    input               PTB_valid_d,            // Valid Data - unregistered
    input               PTB_vc,                 // VC for this packet
    input               PTB_crf,                // CRF for this packet
    input               PTB_in_packet,          // Indicates in packet
    input               PTB_skip_final_crc,     // Indicated to skip final CRC insertion
    input        [15:0] PTB_crc64,              // The current CRC value
    input        [15:0] PTB_crc48,              // The current CRC value
    input        [15:0] PTB_crc32,              // The current CRC value
    input        [15:0] PTB_crc16,              // The current CRC value
    input        [5:0]  PTB_next_fm,            // The ACK ID for this packet
    input               PTB_insert_mid_crc,     // Insert the mid CRC
    input               PTB_mid_crc_inserted,   // A mid CRC was inserted

    // OLLM TX Data Mux Interface
    output reg   [63:0] PTA_data,               // Data
    output reg   [1:0]  PTA_valid_d,            // Early valid indicator
    output reg   [1:0]  PTA_valid,              // Valid Data Present on PTA_data
    output reg          PTA_sop,                // SOP
    output reg          PTA_eop_d,              // Early EOP
    output reg          PTA_eop,                // EOP
    output reg          PTA_in_packet_d,        // Early in a packet indicator
    output reg          PTA_in_packet,          // Currently in a packet

    // OPLM Interface
    input               PP_idle2_selected,      // Indicates the operating idle mode

    // OLLM TX Ready Generator Interface
    output reg          PTA_stall,              // Stall from this module 
    input               PTR_pta_advance         // Advance this module
    // }}} end Port Declarations
  );                  

  // {{{ Local Parameters
  // When in IDLE2 mode, ack id's are 6 bits; for IDLE1 mode only 5 bits
  localparam ID_WIDTH = (IDLE2) ? 6 : 5;
  // }}} end Local Parameters

  // {{{ Wire Declarations
  reg           phy_rst_q = 1;
  reg           insert_crc_stall;   // A stall is needed for the CRC to be appended to a packet
  reg           insert_crc_stall_d; // Inserts a stall in the pipe for the crc to be inserted
  reg           mid_crc_inserted_q;
  // }}} end Wire Declarations

  // {{{ Register Reset
  // Must register the reset before use
  always @(posedge phy_clk) begin
    phy_rst_q <= #TCQ phy_rst;
  end
  // }}} end Register Reset

  // {{{ Stall Generator
  // Generate the stall to pass to the ready generator 
  // 1. We are not stalling to insert an extra cycle for CRC/Pad
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PTA_stall <= #TCQ 0;
    end else begin
      PTA_stall <= #TCQ ((insert_crc_stall_d && PTR_pta_advance && !(PTB_mid_crc_inserted && !PTB_eop)) || 
                         (insert_crc_stall && !PTR_pta_advance));
    end
  end
  // }}} end Ready Generator

  // {{{ Assemble Data w/Valid
  // Prefix the data with the ack id and append on the CRC and optionally PAD
  reg [23:0]  ptb_data_q;
  reg [3:0]   ptb_keep_q;
  reg [15:0]  ptb_crc64_q;
  reg [15:0]  ptb_crc48_q;
  reg [63:0]  pta_data_d;
  reg         pta_in_packet_d;
  reg         pta_sop_d;
  reg         insert_mid_crc_q;

  // Select the first byte dependent on the operating idle mode
  wire [7:0] first_byte = (PP_idle2_selected) ? {PTB_next_fm, PTB_vc, PTB_crf} :
                                                {PTB_next_fm[4:0], 1'b0, PTB_vc, PTB_crf};      

  // Save off the first few bytes to append as needed
  // Only update this for active beats.
  always @(posedge phy_clk) begin
    if (PTB_valid && PTR_pta_advance) begin
      ptb_data_q         <= #TCQ PTB_data[23:0];
      ptb_keep_q         <= #TCQ PTB_keep;
      ptb_crc64_q        <= #TCQ PTB_crc64;
      ptb_crc48_q        <= #TCQ PTB_crc48;
    end
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      mid_crc_inserted_q <= #TCQ 1'b0;
      insert_mid_crc_q   <= #TCQ 1'b0;
    end else if (PTB_valid && PTR_pta_advance) begin
      mid_crc_inserted_q <= #TCQ PTB_mid_crc_inserted;
      insert_mid_crc_q   <= #TCQ PTB_insert_mid_crc;
    end
  end

  // Based on where we are in packet, select the output data
  always @* begin
    PTA_valid_d        = 0;
    pta_sop_d          = 0;
    PTA_eop_d          = 0;
    PTA_in_packet_d    = 0;
    pta_data_d         = 0;
    insert_crc_stall_d = 0;

    casex ({insert_crc_stall, PTB_sop, PTB_eop, PTB_in_packet})
      // Inserted an extra cycle for the mid CRC this will only happen
      // if the strobe was 5 or 7
      // REQ: req_pt_mid_crc16
      // REQ: req_pt_pad_inserted_correctly
      4'b1xxx: begin
        //1 bytes left that is valid
        if (ptb_keep_q[0]) begin
          pta_data_d = (mid_crc_inserted_q || insert_mid_crc_q) ? 
                       {ptb_data_q[23:8], ptb_crc64_q, 32'b0} :
                       {ptb_crc64_q, 48'b0};

        //Just need the crc. If the strobe indicated 5 bytes valid then we
        //need the 48 bit CRC
        // REQ: req_pt_pad_inserted_correctly
        end else begin
          pta_data_d = {ptb_crc48_q, 48'b0};
        end

        PTA_valid_d     = 2'b10;
        PTA_eop_d       = 1;
        PTA_in_packet_d = 1;
      end

      // SOP
      4'b010x: begin
        pta_data_d      = {first_byte, PTB_data[63:8]};
        PTA_valid_d     = {2{PTB_valid}};
        pta_sop_d       = 1;
        PTA_eop_d       = 0;
        PTA_in_packet_d = 1;
      end

      // SOP and EOP
      4'b011x: begin
        //A single cycle packet can only ever have a stobe of 5 or 7 bytes
        //7 Bytes Valid Case
        // REQ: req_pt_end_crc16
        if (PTB_keep[0]) begin 
          pta_data_d         = {first_byte, PTB_data[63:8]};
          insert_crc_stall_d = 1;

        //5 Bytes Valid Case
        end else begin 
          pta_data_d   = {first_byte, PTB_data[63:24], PTB_crc48};
          PTA_eop_d    = 1;
        end
        PTA_valid_d     = {2{PTB_valid}};
        pta_sop_d       = 1;
        PTA_in_packet_d = 1;
      end
       
      // EOP
      4'b001x: begin
        //generate valid and eof based on the strobe
        // REQ: req_pt_end_crc16
        // REQ: req_pt_pad_inserted_correctly
        case (PTB_keep)
          //1 byte is valid
          4'b1000: begin
            PTA_in_packet_d = 1;
            PTA_eop_d       = 1;
            PTA_valid_d     = (PTB_mid_crc_inserted || PTB_insert_mid_crc) ? 
                              2'b11 : 2'b10;

            if (PTB_insert_mid_crc) begin
              pta_data_d   = {ptb_crc64_q, ptb_data_q[7:0], PTB_data[63:56], PTB_crc16,  16'b0};
            end else if (!PTB_mid_crc_inserted) begin
              pta_data_d   = {ptb_data_q[7:0],  PTB_data[63:56], PTB_crc16, 32'b0}; 
            end else begin
              pta_data_d   = {ptb_data_q[23:0], PTB_data[63:56], PTB_crc16, 16'b0};
            end                  
          end
          //3 bytes are valid
          4'b1100: begin
            PTA_in_packet_d = 1;
            PTA_eop_d       = 1;
            PTA_valid_d     = 2'b11;

            if (PTB_insert_mid_crc) begin
              pta_data_d   = {ptb_crc64_q, ptb_data_q[7:0], PTB_data[63:40], PTB_crc32};
            end else if (!PTB_mid_crc_inserted) begin
              pta_data_d   = {ptb_data_q[7:0],  PTB_data[63:40], PTB_crc32, 16'b0}; 
            end else begin
              pta_data_d   = {ptb_data_q[23:0], PTB_data[63:40], PTB_crc32};
            end                   
          end
          //5 bytes are valid
          4'b1110: begin
            PTA_in_packet_d     = 1;
            insert_crc_stall_d = (PTB_mid_crc_inserted || PTB_insert_mid_crc);
            PTA_eop_d          = !(PTB_mid_crc_inserted || PTB_insert_mid_crc); 
            PTA_valid_d        = 2'b11;       

            if (PTB_insert_mid_crc) begin
              pta_data_d   = {ptb_crc64_q, ptb_data_q[7:0], PTB_data[63:24]};
            end else if (!PTB_mid_crc_inserted) begin
              pta_data_d   = {ptb_data_q[7:0],  PTB_data[63:24], PTB_crc48}; 
            end else begin
              pta_data_d   = {ptb_data_q[23:0], PTB_data[63:24]};
            end                      
          end
          //7 bytes are valid
          4'b1111: begin
            PTA_in_packet_d    = 1;
            insert_crc_stall_d = 1;
            PTA_valid_d        = 2'b11;

            if (PTB_insert_mid_crc) begin
              pta_data_d   = {ptb_crc64_q, ptb_data_q[7:0], PTB_data[63:24]};
            end else if (!PTB_mid_crc_inserted) begin
              pta_data_d   = {ptb_data_q[7:0],  PTB_data[63:8]}; 
            end else begin
              pta_data_d   = {ptb_data_q[23:0], PTB_data[63:24]};
            end 
          end

          //Propigate X's for any other strobe value
          default: begin
            PTA_in_packet_d    = 1'bX;
            insert_crc_stall_d = 1'bX;
            PTA_eop_d          = 1'bx;
            PTA_valid_d        = 2'bXX;
            pta_data_d         = 64'hXXXX_XXXX_XXXX_XXXX;
          end
        endcase
      end

      // Mid-pkt
      4'b0001: begin
        // REQ: req_pt_mid_crc16
        if (PTB_insert_mid_crc) begin
          pta_data_d   = {ptb_crc64_q, ptb_data_q[7:0], PTB_data[63:24]};
        end else if (!PTB_mid_crc_inserted) begin
          pta_data_d   = {ptb_data_q[7:0], PTB_data[63:8]};
        end else begin
          pta_data_d   = {ptb_data_q[23:0], PTB_data[63:24]};
        end

        PTA_valid_d     = {2{PTB_valid}};
        PTA_in_packet_d = 1;
      end
    endcase
  end

  //*ASSERTION*
  //(ap_invalid_beat_w_sop): If PTB_sop is asserted valid must also be
  //asserted.
  
  //*ASSERTION*
  //(ap_invalid_beat_w_eop): If PTB_eop is asserted valid must also be
  //asserted.

  //*COVERAGE*
  //(cp_invalid_beat_in_pkt): Cover that an invalid beat is seen in packet

  //*COVERAGE*
  //(cr_pkt_combos): cross all of the following
  //PTB_sop, PTB_eop, PTB_in_packet, insert_crc_stall, ptb_keep_q, PTB_mid_crc_inserted
      
  //*COVERAGE*
  //(cr_midcrc_w_eop): Cross PTB_mid_crc_inserted with eop

  // Register the values
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PTA_valid         <= #TCQ 0;
      PTA_sop           <= #TCQ 0;
      PTA_eop           <= #TCQ 0;
      PTA_in_packet     <= #TCQ 0;
      insert_crc_stall  <= #TCQ 0;

    end else begin
      if (PTR_pta_advance) begin
        PTA_valid         <= #TCQ PTA_valid_d;
        PTA_sop           <= #TCQ pta_sop_d;
        PTA_eop           <= #TCQ PTA_eop_d;
        PTA_in_packet     <= #TCQ PTA_in_packet_d;
        PTA_data          <= #TCQ pta_data_d;
        insert_crc_stall  <= #TCQ insert_crc_stall_d;
      end
    end
  end

  //*ASSERTION*
  //(ap_insert_crc_stall_extended): Insert_crc_stall must only assert for one
  //cycle.

  //*ASSERTION*
  //(ap_insert_crc_stall_inpkt): If insert_crc_stall is asserted then we must
  //be in packet
  // }}} end Assemble Data w/Valid

  // {{{ CRC Check (SWITCH MODE ONLY)
  // Only generate the CRC check if SWITCH MODE was enabled
  generate if (SWITCH_MODE) begin: switch_crc_err_gen
    // Only check the final CRC when:
    // 1. a switch mode core was generated
    // 2. the packet SKIP_CRC bit was asserted indicating
    //    the packet has a final CRC on it.
    reg [15:0] final_crc;

    always @* begin
      case (PTB_keep)
        4'b1000: final_crc = {ptb_data_q[7:0], PTB_data[63:56]};
        4'b1100: final_crc = PTB_data[55:40];
        4'b1110: final_crc = PTB_data[39:24];
        4'b1111: final_crc = PTB_data[23:8];
        default: final_crc = 16'hXXXX;
      endcase
    end

    wire check_crc = PTB_skip_final_crc && PTB_eop;
    wire crc_error = (final_crc != PTB_crc64);

    always @(posedge phy_clk) begin
      if (phy_rst_q) begin
        PT_switch_crc_err <= #TCQ 0;
      end else begin
        if (check_crc && crc_error) begin
          PT_switch_crc_err <= #TCQ 1;
        end else begin
          PT_switch_crc_err <= #TCQ 0;
        end
      end
    end

  // Drive this to 0 if SWITCH MODE is not supported
  end else begin: no_switch_crc_err_gen
    always @(posedge phy_clk) begin
      PT_switch_crc_err <= #TCQ 0;
    end
  end endgenerate //end if (SWITCH_MODE)

  //*COVERAGE*
  // (cp_all_strobes_w_switchmode): Cover al the expected strobes when switch mode is enabled    
  // }}} end CRC Check
endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/phy/ollm_tx/srio_gen2_v4_1_16_ollm_tx_oplm.v#1 $
//----------------------------------------------------------------------
//
// OLLM_TX_OPLM
// Description:
// This module interface with the oplm to provided the appropriate 
// handshaking for link requests and clock compensation
//
// Hierarchy:
// PHY_TOP
//    |___OLLM_TX_TOP
//             |_____OLLM_TX_READY_GEN
//             |_____OLLM_TX_BUF
//             |_____OLLM_TX_PKT_ASSEMBLY
//             |_____OLLM_TX_CS_GEN
//             |_____OLLM_TX_DATA_MUX
//             |_____OLLM_TX_OPLM  <-- this module
// ---------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_ollm_tx_oplm
  #(
    parameter TCQ         = 100 
  )
  (
    // {{{ Port Declarations
    // System Signals
    input               phy_clk,              // PHY interface clock
    input               phy_rst,              // Reset for PHY clock Domain

    // OLLM TX Data Mux Interface
    input       [63:0]  PTM_data,             // Data
    input       [1:0]   PTM_valid,            // Data Valid
    input       [7:0]   PTM_charisk,          // K character locations in Data
    input               PTM_send_lreq,        // Data is a link request

    // OPLM TX Interface Signals
    output reg  [63:0]  PTP_tx_data,          // Transmit data
    output reg  [7:0]   PTP_tx_charisk,       // Indicates which bytes  are K characters
    output reg  [1:0]   PTP_tx_valid,         // Indicates valid words
    input               PP_ccomp_req,         // Request break for clock compensation sequence
    output reg          PTP_ccomp_grant,      // Insert clock compensation at next invalid
    output reg          PTP_send_lreq,        // Indicates the data on PT_tx_data is a LREQ
    input               PP_lreq_sent,         // Indicates the LREQ SYNC SEQ was sent

    // OLLM TX Ready Generator Interface
    output reg          PTP_stall,            // Stall Indicator from this module
    input               PTR_ptp_advance       // Advance this module
    // }}} end Port Declarations
  );                  
  
  // {{{ Wire Declarations
  reg   phy_rst_q = 1;

  reg   pp_lreq_sent_q;   // Registered version on pp_lreq_sent
  reg   lreq_stall;       // A stall is required for a link request to be held
  reg   lreq_stall_q;     // Registered version of lreq_stall
  reg   ccomp_grant_d;    // Insert a stall for the ccomp sequence
  // }}} end Wire Declarstion

  // {{{ Register Reset
  // Must register the reset before use
  always @(posedge phy_clk) begin
    phy_rst_q <= #TCQ phy_rst;
  end
  // }}} end Register Reset

  // {{{ LREQ Stall Generation
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      pp_lreq_sent_q <= #TCQ 0;
    end else begin
      pp_lreq_sent_q <= #TCQ PP_lreq_sent;
    end
  end

  // Stall for a link request as soon as it arrives and hold it until
  // the OPLM indicates it was sent by deasserting the PP_lreq_sent signal
  always @* begin
    if (!pp_lreq_sent_q && PP_lreq_sent) begin
      lreq_stall = 0;

    end else if (PTM_send_lreq && PTR_ptp_advance) begin
      lreq_stall = 1;

    end else begin
      lreq_stall = lreq_stall_q;
    end
  end

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      lreq_stall_q <= #TCQ 0;
    end else begin
      lreq_stall_q <= #TCQ lreq_stall;
    end
  end
  // }}} end LREQ Stall Generation

  // {{{ CCOMP Grant Generation
  // Grant clock compensation insertion when it has been requested and there
  // is gap in the data.
  always @* begin
    if (!PP_ccomp_req) begin
      ccomp_grant_d = 1'b0;

    //When there is a gap in valid data arriving and any current data was
    //already accepted, assert the grant for the ccomp sequence
    end else if (PP_ccomp_req && !(|PTM_valid) && !(|PTP_tx_valid)) begin
      ccomp_grant_d = 1'b1;
    
    end else begin
      ccomp_grant_d = PTP_ccomp_grant;
    end
  end

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PTP_ccomp_grant <= #TCQ 0;
    end else begin
      PTP_ccomp_grant <= #TCQ ccomp_grant_d;
    end
  end
  // }}} end CCOMP Grant Generation

  // {{{ Stall Generation
  // This module stalls for:
  // 1. LREQ tranmission
  // 2. CCOMP_REQ assertion
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PTP_stall <= #TCQ 0;
    end else begin
      PTP_stall <= #TCQ lreq_stall || ccomp_grant_d;
    end
  end
  // }}} end Ready Generation

  // {{{ Register Outputs
  //Drive Data to the OPLM TX Interface
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PTP_tx_valid    <= #TCQ 0;
      PTP_send_lreq   <= #TCQ 0;
    end else begin
      if (!lreq_stall && lreq_stall_q) begin
        PTP_tx_valid    <= #TCQ 2'b0;
        PTP_send_lreq   <= #TCQ 1'b0;

      end else if (PTR_ptp_advance) begin
        PTP_tx_data     <= #TCQ PTM_data;
        PTP_tx_charisk  <= #TCQ PTM_charisk;
        PTP_tx_valid    <= #TCQ PTM_valid;
        PTP_send_lreq   <= #TCQ PTM_send_lreq;
      end
    end
  end
  // }}} Register Outputs

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/phy/ollm_tx/srio_gen2_v4_1_16_ollm_tx_data_mux.v#1 $
//----------------------------------------------------------------------
//
// OLLM_TX_DATA_MUX
// Description:
// This module is responsible for accepting the packets from  
// packet assembly and control symbol generation and muxing them into
// one complete data stream with no gaps in between when possible.
//
// Hierarchy:
// PHY_TOP
//    |___OLLM_TX_TOP
//             |_____OLLM_TX_READY_GEN
//             |_____OLLM_TX_BUF
//             |_____OLLM_TX_PKT_ASSEMBLY
//             |_____OLLM_TX_CS_GEN 
//             |_____OLLM_TX_DATA_MUX <-- this module
//             |_____OLLM_TX_OPLM
// ---------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_ollm_tx_data_mux
  #(
    parameter TCQ = 100 
  )
  (
    // {{{ Port Declarations
    // System Signals
    input               phy_clk,            // PHY interface clock
    input               phy_rst,            // Reset for PHY clock Domain

    // Inputs required for bind file
    input               PT_phy_rewind,      // A rewind is in progress
    
    // OLLM TX Data Mux Interface
    input        [63:0] PTA_data,           // Data
    input        [1:0]  PTA_valid_d,        // Early valid
    input        [1:0]  PTA_valid,          // Valid Data Present on PTB_data
    input               PTA_sop,            // SOP
    input               PTA_in_packet_d,    // Early In Packet
    input               PTA_in_packet,      // In Packet
    input               PTA_eop_d,          // Early EOP
    input               PTA_eop,            // EOP

    // OLLM TX CS Gen Interface
    input        [63:0] PTS_data,           // Data
    input        [1:0]  PTS_valid,          // Valid Data Present on PTB_data
    input               PTS_lreq,           // Indicates the data is a link request
    input               PTS_embed_cs,       // Indicates to send the control symbol immediately
    input        [7:0]  PTS_charisk,        // Indicates which bytes are K characters
    input               PTS_sop,            // Indicates an SOP 
    input               PTS_eop,            // Indicates an EOP 

    // OLLM RX Interface
    input               PR_link_initialized,// Link is Init, needed for bind file 

    // OPLM Interface
    output reg   [1:0]  PTM_tx_early_valid, // Early valid indicator for the OPLM
    output reg          PTM_tx_early_lreq,  // Early lreq indicator for the OPLM
    input               PP_ccomp_req,       // Indicates a Clk Comp. Sequence is needed  
    input               PP_idle2_selected,  // Operating Idle mode

    // OLLM TX OPLM Interface
    output reg   [63:0] PTM_data,           // Data
    output reg   [1:0]  PTM_valid,          // Data Valid
    output reg   [7:0]  PTM_charisk,        // K character locations in Data
    output reg          PTM_send_lreq,      // Data is a link request

    // OLLM TX Ready Generator Interface
    output reg          PTM_pta_stall,      // Stall the Packet Data
    output reg          PTM_pts_stall,      // Stall the Control Symbol Generator
    input               PTR_pta_advance,    // Advance the Packet Assembly
    input               PTR_pts_advance,    // Advance the Control Symbol Generator
    input               PTR_ptm_advance     // Advance the Data Mux
    // }}} end Port Declarations
  );     

  // {{{ Local Parameters
  // Local params used to select the data output of this module 
  // from packet assembly and the control symbol generator.
  localparam PTS_PTS = 2'b00;   // All CSG data
  localparam PTS_PTA = 2'b01;   // First half CSG data, second half PAM data
  localparam PTA_PTS = 2'b10;   // First half PAM data, second half CSG Data
  localparam PTA_PTA = 2'b11;   // All PAM data
  // }}} end Local Parameters
 
  // {{{ Wire Declarations
  reg           phy_rst_q = 1;

  // The half of the packet data which was accepted but not sent yet
  reg   [31:0]  pta_data_q;
  reg           pta_eop_q;
  reg           pta_active_q;
  reg           pta_shifted;
  wire          pta_eop_active;
  wire          pta_dead_beat_d;
  reg           pta_dead_beat;
  reg           pta_dead_beat_q;
  reg           pta_dead_beat_qq;

  // The half of the control symbol data which was accepted but not yet sent.
  reg   [31:0]  pts_data_q;
  reg           pts_valid_q;
  reg   [3:0]   pts_charisk_q;
  reg           pts_shifted;
  reg           pts_sop_q;

  // Packet Data shifting signals
  wire [63:0]   pta_data_realigned;
  wire          pta_valid_lower_bit;
  reg  [1:0]    pta_valid_realigned;

  // No K characters in packets
  wire [7:0]    pta_charisk_realigned;
  

  // Control symbol shifting signals
  reg   [1:0]   pts_valid_realigned;
  wire          pts_embed_active;
  wire          accept_embed_cs;
  reg           accept_embed_cs_q;
  wire  [63:0]  pts_data_realigned;
  wire  [7:0]   pts_charisk_realigned;

  // The shifted version of the data to transmit
  reg   [63:0]  data_realigned;
  reg   [1:0]   valid_realigned;
  reg   [7:0]   charisk_realigned; 

  // Control signals for in packet scenarios 
  reg   [1:0]   oopkt_data_select;
  reg           oopkt_pta_shifted_d;
  reg           oopkt_pts_shifted_d;
  reg           oopkt_pts_stall_d;
  reg           oopkt_pta_stall_d;

  // Control signals for out of packet scenarios
  reg   [1:0]   inpkt_data_select;
  reg           inpkt_pta_shifted_d;
  reg           inpkt_pts_shifted_d;
  reg           inpkt_pts_stall_d;
  reg           inpkt_pta_stall_d;

  wire  [1:0]   data_select;        // What kind of data to select
  reg           in_packet_sel;      // In packet select
  wire  [1:0]   pta_active;         // Active PTA cycle
  reg           pta_ccomp_stall;    // Stall packet data for the ccomp seq
  reg           pta_ccomp_stall_q;  // registered pta_ccomp_stall
  reg           pts_ccomp_stall;    // Stall control symbols for the ccomp seq
  reg           pts_ccomp_stall_q;  // registered pts_ccomp_stall
  reg           ccomp_req_q_advance;// ccomp stall value only on advance
  wire          ccomp_req_rose;     // rising edge of ccomp stall for active cycles
  // }}} end Wire Declarations

  // {{{ if SIMULATION
  // Make data selection types readable in the waveform for
  // simulation/debugging
  `ifdef SIMULATION
    reg [15*8-1:0] data_select_string = "null";

    always @* begin
      //Data Select Decode
      case (data_select)
        PTS_PTS: data_select_string = "PTS_PTS";
        PTS_PTA: data_select_string = "PTS_PTA";
        PTA_PTS: data_select_string = "PTA_PTS";
        PTA_PTA: data_select_string = "PTA_PTA";
        default: data_select_string = "INVALID";
      endcase
    end
  `endif
  // }}} end if SIMULATION

  // {{{ Register Reset
  // Must register the reset before use
  always @(posedge phy_clk) begin
    phy_rst_q <= #TCQ phy_rst;
  end
  // }}} end Register Reset

  // {{{ Clock Compensation Stalling Logic
  // Figure out when to mask off transmitting when a clock compensation needs
  // to be inserted.

  // Start stalling once the EOP has been inserted if we were in packets,
  // Otherwise start stalling if there is no valid data pending.
  assign ccomp_req_rose = PP_ccomp_req && !ccomp_req_q_advance;

  always @* begin
    if (!PP_ccomp_req || (PTR_pts_advance && PTS_sop)) begin
      pta_ccomp_stall =  0;
    end else if (((PTA_valid == 2'b00 && PTS_valid == 2'b00 && !PTA_in_packet) || 
                  (PTA_eop && PTR_pta_advance && !PTS_sop && !ccomp_req_rose) ||
                  (PTS_eop && PTR_pts_advance)) && PP_ccomp_req) begin
      pta_ccomp_stall = 1;
    end else begin
      pta_ccomp_stall = pta_ccomp_stall_q;
    end
  end

  always @* begin
    if (!PP_ccomp_req) begin
      pts_ccomp_stall =  0;
    end else if (((PTA_valid == 2'b00 && PTS_valid == 2'b00 && !PTA_in_packet) || 
                  (PTS_eop && PTR_pts_advance)) && PP_ccomp_req) begin
      pts_ccomp_stall = 1;
    end else begin
      pts_ccomp_stall = pts_ccomp_stall_q;
    end
  end
  
  // Latch the ccomp stall signal
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      pta_ccomp_stall_q   <= #TCQ 0;
      pts_ccomp_stall_q   <= #TCQ 0;
      ccomp_req_q_advance <= #TCQ 0;
    end else begin
      pta_ccomp_stall_q <= #TCQ pta_ccomp_stall;
      pts_ccomp_stall_q <= #TCQ pts_ccomp_stall;

      // Only sample when advancing to look for the rising edge
      if (PTR_pta_advance)
        ccomp_req_q_advance  <= #TCQ PP_ccomp_req;
    end
  end

    
  //*COVERAGE*
  //(cp_pta_before_pts_ccomp_stall): See a ccomp stall on the packet data before the
  // control symbol data

  //*COVERAGE*
  //(cp_pta_pts_ccomp_stall): See a ccomp stall on both the packet data and the
  // control symbol data

  //*ASSERTION*
  //(ap_pts_before_pta_ccomp_stall): There should never be a control symbol stall
  // before a data stall

  // }}} end Clock Compensation Stalling Logic

  // {{{ PAM/CSG Data Shifting
  // Save off the lower half of the data from Packet Assembly in case it 
  // needs to be shifted 
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      pta_eop_q    <= #TCQ 0;
      pta_data_q   <= #TCQ 0;
      pta_active_q <= #TCQ 0;
    end else begin
      if (PTR_pta_advance) begin
        pta_eop_q    <= #TCQ PTA_eop;
        pta_data_q   <= #TCQ PTA_data[31:0];
        pta_active_q <= #TCQ PTA_valid[0];
      end
    end
  end

  // Shift the data from PAM as needed
  assign pta_active            = {PTA_valid[1] & PTR_pta_advance, 
                                  PTA_valid[0] & PTR_pta_advance};
  assign pta_data_realigned    = (pta_shifted) ? {pta_data_q,  PTA_data[63:32]} : PTA_data;

  // Mask off the lower bits valid if the data is shifted and we are starting a new packet
  assign pta_valid_lower_bit   = (PTA_sop) ? 0 : PTA_valid[1] || 
                                                 (pta_shifted && PTA_eop && PTA_valid[1]);

  always @* begin
    if (pta_shifted && pta_dead_beat_qq) begin
      pta_valid_realigned = {1'b1, pta_valid_lower_bit};
    end else if (pta_shifted) begin
      pta_valid_realigned = {pta_active_q, pta_valid_lower_bit};
    end else begin
      pta_valid_realigned = PTA_valid;
    end
  end

  // No K characters in packets
  assign pta_charisk_realigned = 8'b0;

  // Save off the lower half of the data from the Control Symbol Generator
  // in case it needs to be shifted.
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      pts_data_q    <= #TCQ 0;
      pts_valid_q   <= #TCQ 0;
      pts_charisk_q <= #TCQ 0;
      pts_sop_q     <= #TCQ 0;
    end else begin
      pts_data_q    <= #TCQ PTS_data[31:0];
      pts_valid_q   <= #TCQ PTS_valid[0];
      pts_charisk_q <= #TCQ PTS_charisk[3:0];
      pts_sop_q     <= #TCQ PTS_sop;
    end
  end

  // Shift the data from CSG as needed
  assign pts_data_realigned    = (pts_shifted) ? {pts_data_q,   PTS_data[63:32]} : PTS_data;
  assign pts_charisk_realigned = (pts_shifted) ? {pts_charisk_q,PTS_charisk[7:4]}: PTS_charisk;
  assign accept_embed_cs       = PTS_embed_cs && !(PTS_sop || PTS_eop) && !PTR_pts_advance;
  assign pts_embed_active      = accept_embed_cs_q && PTR_pts_advance;
  wire   pts_valid_lower_bit   = (pts_sop_q || (pts_ccomp_stall_q && !PTS_eop) || 
                                  (!PTR_pts_advance && pts_shifted)) ? 
                                    0 :  PTS_valid[1];


  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      accept_embed_cs_q <= #TCQ 0;
    end else begin
      accept_embed_cs_q <= #TCQ accept_embed_cs;
    end
  end

  always @* begin
    // Wait until after an EOP before masking the control symbols to be sure
    // a packets complete before starting the ccomp sequence
    if (pts_ccomp_stall_q && !PTS_eop && !pts_shifted) begin
      pts_valid_realigned = 0;

    end else if (PTA_in_packet && !PTA_eop && !(|PTA_valid)) begin
      pts_valid_realigned = (pta_shifted && !PP_idle2_selected) ? 2'b10 : 2'b11;
    
    // If a dead beat was inserted, it will only be shifted for a full dword
    // of control symbols, if this is the case make the upper bit valid for
    // the second half of the dword
    end else if (pts_shifted && pta_dead_beat_q) begin
      pts_valid_realigned = {1'b1,  pts_valid_lower_bit};

    end else begin
      pts_valid_realigned = (pts_shifted) ? {pts_valid_q,  pts_valid_lower_bit} : PTS_valid;
    end
  end

  // Check for an active EOP so we know when to move out of packet. need to
  // account for the end of an arriving packet which was shifted and if a dead
  // beat was inserted directly before the EOP
  assign pta_eop_active = (pta_shifted && &PTA_valid) ? pta_eop_q && PTR_ptm_advance : 
                                                        PTA_eop && PTR_pta_advance && 
                                                          !(pts_embed_active && &PTA_valid) &&
                                                          !(&PTA_valid && pts_shifted && pta_dead_beat_q);

  // Logic to toggle between in packet and out of packet selection.
  // Needs to account for two half dwords for single cycle packets.
  wire tiny_pkt_toggle = (PTA_eop && PTA_sop && |pta_active) && 
                         !(^pts_valid_realigned && ^pta_valid_realigned);

  wire ending_pkt_toggle = ((pta_eop_active && 
                            !(^pts_valid_realigned && ^pta_valid_realigned && PTS_sop && PTR_pts_advance)) || 
                            !PTA_in_packet);

  // Move into packet if we accept an SOP
  // This will be PTS_sop being accepted in the case where the control symbol
  // is aligned. This will be PTA_sop being accepted in the case where the
  // control symbol was shifted and now we started accepting data.
  wire starting_pkt_toggle = (PTS_sop && PTR_pts_advance && (!pts_shifted || !(&PTS_valid))) || 
                             (PTA_sop && PTR_pta_advance && pts_shifted);

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      in_packet_sel <= #TCQ 0;
    end else begin
      if (PTR_ptm_advance) begin
        if (pta_ccomp_stall && pts_ccomp_stall) begin
          in_packet_sel <= #TCQ 0;

        end else if (tiny_pkt_toggle) begin
          in_packet_sel <= #TCQ ~in_packet_sel;

        end else if (ending_pkt_toggle && in_packet_sel) begin
          in_packet_sel <= #TCQ 0;

        end else if (starting_pkt_toggle && !in_packet_sel) begin
          in_packet_sel <= #TCQ 1;
        end
      end //end if (PTR_ptm_advance)
    end
  end

  // Based on the Data Select signal, mux the control symbol with the packet
  // to form the new stream.
  assign data_select = (in_packet_sel) ? inpkt_data_select : oopkt_data_select;

  always @* begin
    case (data_select)
      PTS_PTS: begin
        data_realigned    = pts_data_realigned;
        valid_realigned   = pts_valid_realigned;
        charisk_realigned = pts_charisk_realigned;
      end

      PTS_PTA: begin
        data_realigned    = {pts_data_realigned[63:32], pta_data_realigned[63:32]};
        valid_realigned   = {pts_valid_realigned[1],    pta_valid_realigned[1]};
        charisk_realigned = {pts_charisk_realigned[7:4],pta_charisk_realigned[7:4]};
      end

      PTA_PTS: begin
        data_realigned    = {pta_data_realigned[63:32], pts_data_realigned[63:32]};
        valid_realigned   = {pta_valid_realigned[1],    pts_valid_realigned[1]};
        charisk_realigned = {pta_charisk_realigned[7:4],pts_charisk_realigned[7:4]};
      end

      PTA_PTA: begin
        data_realigned    = pta_data_realigned;
        valid_realigned   = pta_valid_realigned;
        charisk_realigned = pta_charisk_realigned;
      end

      default: begin
        data_realigned    = {64{1'bX}};
        valid_realigned   = {2{1'bX}};
        charisk_realigned = {8{1'bX}};
      end
    endcase
  end  
  
  //*ASSERTION*
  //(cp_cs_inserted_wo_advance0/cp_cs_inserted_wo_advance1): If a valid control symbol is 
  // inserted into the data stream, PTR_pts_advance must be asserted

  //*ASSERTION*
  //(ap_pts_advance_in_packet): If a control symbol is accepted then the data
  //mux must be currently accepting it.

  //*COVERAGE*
  //(cr_data_select): Cover all cases of data selection and the pts_shifted
  //and pta_shifted control signals with embedding control symbols
  

  // Indicate when an in packet dead beat is arriving
  assign pta_dead_beat_d = (PTA_valid_d == 2'b00) && PTA_in_packet_d && PTR_pta_advance;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      pta_dead_beat    <= #TCQ 0;
      pta_dead_beat_q  <= #TCQ 0;
      pta_dead_beat_qq <= #TCQ 0;
    end else begin
      pta_dead_beat    <= #TCQ pta_dead_beat_d;
      pta_dead_beat_q  <= #TCQ pta_dead_beat;
      pta_dead_beat_qq <= #TCQ pta_dead_beat_q;
    end
  end

  //*COVERAGE*
  //(cp_dead_beat_idle1): Observe a dead beat in idle1 

  //*COVERAGE*
  //(cp_dead_beat_idle1): Observe a dead beat in idle2

  //*COVERAGE*
  //(cp_b2b_dead_beats_idle1): See back to back dead beats in idle1

  //*COVERAGE*
  //(cp_b2b_dead_beats_idle2): See back to back dead beats in idle2

  //*COVERAGE*
  //(cp_dead_beat_before_eop): See a beat beat followed by EOP

  //*COVERAGE*
  //(cp_dead_beat_after_sop): See a beat beat follow SOP

  //*COVERAGE*
  //(cp_dead_beat_w_embed_cs_idle1): See a dead beat occur with an embeded control symbol in idle1

  //*COVERAGE*
  //(cp_dead_beat_w_embed_cs_idle2): See a dead beat occur with an embeded control symbol in idle2

  // }}} end PAM/CSG Data Shifting
  
  // {{{ + Data Mux Control Logic +
  
  // {{{ Out of Packet Select
 // Calculate the next values for the out of packet scenarios
  always @* begin
    oopkt_pta_shifted_d = pta_shifted;
    oopkt_pts_shifted_d = pts_shifted;
    oopkt_pts_stall_d   = 0;
    oopkt_pta_stall_d   = 0;

    casex ({PTS_lreq, pts_valid_realigned})
      // If there is a shifted link-request we need to unshift before sending
      3'b1_XX: begin
        oopkt_data_select   = PTS_PTS;
        oopkt_pts_shifted_d = 0;
        oopkt_pta_shifted_d = 0;
        oopkt_pts_stall_d   = pta_ccomp_stall;
      end

      // If only one is valid control symbol set, the data must follow on bits [31:0],
      // if any exists.  Indicate a data shift if we about to be in_packet.
      // Continue to be ready to accept control symbols we are not going to be
      // in packet
      3'b0_10: begin
        // Only select control symbols if we need to start holding off data for
        // the ccomp sequence
        oopkt_data_select   = (pta_ccomp_stall_q || !PTR_pta_advance) ? PTS_PTS : PTS_PTA;
        oopkt_pts_shifted_d = 0;

        // Only shift the packet data if there is valid data which will begin
        // shifting
        oopkt_pta_shifted_d = PTA_valid[1] && !pta_ccomp_stall_q && PTR_pta_advance;

        // Only stall control symbols if we are going in packet and this symbol
        // was accepted, or if the clk compensation sequence was requested.
        // Do not stall if the next in packet cycle there is not valid data.
        oopkt_pts_stall_d   = pts_ccomp_stall || 
                              ((!PTA_eop && PTA_valid[1] && PTR_pta_advance) && !pta_dead_beat_d);

        // Stall packet data if this is the end of the packet if:
        // 1. there is a really small packet
        // 2. to insert the clock compensation sequence
        // 3. packet sop and cs sop are stalled.
        oopkt_pta_stall_d = (PTA_eop && PTR_pta_advance) || pta_ccomp_stall || 
                            (&PTS_valid && !PTR_pts_advance && !PTR_pta_advance);
      end

      // In either case of no valid control symbols or only valid control
      // symbols, always select them
      default: begin
        oopkt_data_select   = PTS_PTS;
        oopkt_pta_shifted_d = 0;

        // The last part stalls in idle2 after EOPs to line up oopkt data in case an LREQ follows
        // the EOP
        oopkt_pts_stall_d   = pts_ccomp_stall || 
                              (PTS_sop && PTR_ptm_advance) || 
                              (pts_shifted && PTS_eop && PTR_pts_advance && PP_idle2_selected);


        oopkt_pta_stall_d   = pta_ccomp_stall || 
                              (|PTA_valid && !PTS_sop && PTR_pts_advance) ||
                              (!PTR_ptm_advance && &PTS_valid) ||
                              (PTA_valid[1] && !PTS_sop);

        //Unshift the control symbols when 
        // 1. there is no valid cs's sitting here
        // 2. we are ending a packet we need to unshift in case an LREQ needs
        //    to be send which needs to be aligned for IDLE2 mode
        if (pts_shifted && (!PTS_valid[0] || PTS_lreq))
          oopkt_pts_shifted_d = 0;
        else
          oopkt_pts_shifted_d = pts_shifted;
      end
    endcase
  end 

  //*COVERAGE*
  //(cp_single_cycle_pkt_start_stall_idle2): Cover a single cycle pkt is seen when the data mux is
  // out of packet and a control symbol is valid that is not the start of the packet in IDLE2

  //*COVERAGE*
  //(cp_single_cycle_pkt_start_stall_idle1): Cover a single cycle pkt is seen when the data mux is
  // out of packet and a control symbol is valid that is not the start of the packet in IDLE1

  // }}} end Out of packet Select
 
  // {{{ In Packet Select
  // Calculate the next values for in packet scenarios
  always @* begin
    inpkt_pta_shifted_d = pta_shifted;
    inpkt_pts_shifted_d = pts_shifted;
    inpkt_pta_stall_d   = 0;
    inpkt_pts_stall_d   = 0;

    casex ({pta_valid_realigned, pts_embed_active, pts_valid_realigned})
      // Full Cycle of Valid Data 
      5'b11_0_XX: begin
        // If the control symbols shifted then full dword of cs was inserted
        // for a dead beat. in this case we need to insert the second half
        inpkt_data_select   = (pts_shifted && pta_dead_beat_q) ? PTS_PTA : PTA_PTA;
        inpkt_pta_shifted_d = (pts_shifted && pta_dead_beat_q) ? 1 : 
                                (pta_eop_active) ? 0 : pta_shifted;
        inpkt_pts_shifted_d = 0;

        // If this was a shifted active last beat, unshift the data going before 
        // going out of packet. Stall packets if we are stating the clock comp sequence
        // or it will take a whole cycle to insert control symbols when we are
        // out of packet.
        if (pta_eop_active) begin
          //inpkt_pta_shifted_d = 0;
          inpkt_pta_stall_d = (PP_ccomp_req && !PTS_sop) || &PTS_valid || PP_idle2_selected;
        
        // Stall packets if we are about to accept embedding a control symbol
        // or EOP is inactive meaning the data was shifted and we need an
        // extra cycle to complete.
        end else begin
          // Stall PTA if:
          // 1. We are accepting an embededd control symbol to be inserted on the next cycle
          // 2. A one-dword EOP is on the next cycle and the CS will be inserted with it
          // 4. Next cycle the EOP will be accepted.
          // 5. A clock compensation needs to be inserted
          inpkt_pta_stall_d = (accept_embed_cs && !pta_dead_beat_d && PTR_pta_advance &&
                                (((PP_idle2_selected || &PTS_valid) && 
                                  !(PTA_eop_d && PTA_valid_d == 2'b10) && PTR_pta_advance) || 
                                 pta_shifted)) ||
                              (PTA_eop && PTR_pta_advance) ||
                              pta_ccomp_stall;
        
          // Do not stall control symbols if:
          // 1. We are going to accept an embedded control symbol
          // 2. On the next cycle is EOP and we need to start the oop control symbols
          // 3. On the next cycle is a dead in packet beat so we need to fill
          //    it with a control symbol
          inpkt_pts_stall_d = !(accept_embed_cs ||
                                (PTA_eop_d && !(&PTA_valid_d) && !pta_shifted && !(pts_shifted && pta_dead_beat_q)) ||
                                (PTA_eop && pta_shifted) ||
                                (pta_dead_beat_d) ||
                               (pts_shifted && pta_dead_beat_q) && PTA_eop) ||
                               !PTR_ptm_advance;
        end
      end

      // Valid data with a long control symbol/two short control symbols
      // that need to be embedded
      5'b11_1_11: begin
        inpkt_data_select = PTS_PTS;
        // Stall control symbol unless the next beat is an in pkt dead beat.
        inpkt_pts_stall_d = !pta_dead_beat_d;
      end

      // Valid data with a short control symbol to embed.
      // If the data was not shifted, it now needs to be shifted.
      // If the data was already shifted, it can now be unshifted.
      // A stall on packet data is needed to insert the control symbol only if
      // not yet shifted. 
      5'b11_1_10: begin
        inpkt_data_select   = PTA_PTS;
        inpkt_pta_shifted_d = ~pta_shifted;
        inpkt_pts_stall_d   = !((PTA_eop && !PTR_pta_advance && !(&PTA_valid)) || 
                                (PTA_eop && PTR_pta_advance && !pta_shifted) || 
                                pta_dead_beat_d);
        inpkt_pta_stall_d   = PTA_eop && PTR_pta_advance;
      end

      // This is either EOP with a short EOP control symbol, or a shifted invalid 
      // data beat which will need to be padded with a short control symbol.
      // In either case, unshift the data and insert the control symbol.
      5'b10_X_10: begin
        inpkt_data_select   = (pts_shifted && pta_dead_beat_q) ? PTS_PTA : PTA_PTS;
        inpkt_pts_shifted_d = (pts_shifted && pta_dead_beat_q) ? 0       : pts_shifted;
        inpkt_pta_shifted_d = (pts_shifted && pta_dead_beat_q && !pta_eop_active);

        //Stall packet data directly following eop if a clock comp is
        //requested, or if we need to insert SOP on the next cycle
        inpkt_pta_stall_d = (pta_ccomp_stall && pta_eop_active) || !PTR_ptm_advance || 
                            (!PTR_pts_advance && &PTS_valid);

        // Stall the cs if:
        // 1. If sop is inserted meaning we are starting in packet
        // 2. This was an in_packet_dead beat and the next cycle is valid, but
        //    only if the next cycle is not a dword size eop.
        // 3. If the clk compensation must be inserted 
        inpkt_pts_stall_d = (PTS_sop && PTR_pts_advance) ||
                            (pta_dead_beat && !pta_dead_beat_d && !(PTA_eop_d && !(&PTA_valid_d))) ||
                            pts_ccomp_stall;
      end

      // This is either EOP with a long EOP control symbol, or a shifted invalid 
      // data beat which will need to be padded with a control symbol.
      // In either case, unshift the data and insert the control symbol. 
      5'b10_X_11: begin
        inpkt_data_select   = (pts_shifted && pta_dead_beat_q) ? PTS_PTA : PTA_PTS;
        inpkt_pta_shifted_d = 0;

        //Stall packet data directly following eop if a clock comp is
        //requested. 
        inpkt_pta_stall_d = pta_ccomp_stall || (!(PTS_sop || PTS_eop) && !pta_dead_beat);

        // Stall the cs if:
        // 1. If sop is inserted meaning we are starting in packet
        // 2. This was an in_packet_dead beat and the next cycle is valid
        // 3. We are sending ending a pkt with a long control symbol.
        //    we need to unshifted cs's so lreqs will always be aligned
        // 4. If the clk compensation must be inserted
        inpkt_pts_stall_d = (PTS_sop && PTR_pts_advance) || 
                            (pta_dead_beat && !pta_dead_beat_d) ||
                            (PP_idle2_selected && PTS_eop) || 
                            pts_ccomp_stall;

        inpkt_pts_shifted_d = 1;
      end

      // Data's EOP ended on the last cycle OR there was a gap in the
      // packet, which was not detectable by the in_packet logic. Insert a
      // control symbol in this case. If were are in packet then there will
      // be a status symbol which will be a filler for the data.
      5'b00_X_XX: begin
        inpkt_data_select   = PTS_PTS;
        inpkt_pta_shifted_d = 0;

        // Stall control symbols if we are still in packet and the next beat
        // is valid and its not going to be an EOP which needs half a control
        // symbol
        inpkt_pts_stall_d = (pta_dead_beat && !pta_dead_beat_d) && 
                            (!(PTA_eop_d && PTA_valid_d == 2'b10) || pts_shifted);
      end

      // Any other case is invalid and X's should be propigated.
      default: begin
        inpkt_data_select   = {2{1'bX}};
        inpkt_pta_shifted_d = 1'bX;
        inpkt_pts_shifted_d = 1'bX;
        inpkt_pts_stall_d   = 1'bX;
        inpkt_pta_stall_d   = 1'bX;
      end
    endcase
  end

  //*COVERAGE*
  //(cr_embed_X_ccomp): cross accepting an embedded control symbol with the
  //clock comp sequence request.

  //*COVERAGE*
  //(cp_embed_two_short): Cover the case where two short control symbols need
  //to be embedded in a packet.

  //*COVERAGE*
  //(cp_embed_one_long): Cover the case where one long control symbol needs to
  //be embedded in a packet

  //*ASSERTION*
  // (ap_embedded_sop_rcvd): An SOP can not be embedded in a packet

  //*ASSERTION*
  // (ap_rewind_without_packet_delimiter): If a rewind occurs in packet, then
  // there must be a control symbol available to kill the packet with.
  // }}} end In Packet Select

  // Register the control signals for this module based on being in a packet
  // or out of packet
  // REQ: req_pt_no_cs_before_port_init

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      pta_shifted <= #TCQ 0;
      pts_shifted <= #TCQ 0;
    end else begin
      if (PTR_ptm_advance) begin
        pta_shifted <= #TCQ (in_packet_sel) ? inpkt_pta_shifted_d : oopkt_pta_shifted_d;
        pts_shifted <= #TCQ (in_packet_sel) ? inpkt_pts_shifted_d : oopkt_pts_shifted_d;
      end
    end
  end 

  // Drive the stalls's back to the ready generator. These are register in the
  // advance signal indicator to the other modules
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PTM_pts_stall <= #TCQ 0;
      PTM_pta_stall <= #TCQ 0;
    end else begin
      PTM_pts_stall <= #TCQ (in_packet_sel) ? inpkt_pts_stall_d : oopkt_pts_stall_d;
      PTM_pta_stall <= #TCQ (in_packet_sel) ? inpkt_pta_stall_d : oopkt_pta_stall_d;
    end
  end

  //*ASSERTION*
  //(ap_pts_shifted_inpkt): pts_shifted should never be true while in packet.

  //*COVERAGE*
  //(cr_input_valid_combos): Cover all combinations of inputs of the valid signals
  //from packet assembly and control symbol generation
   
  //*COVERAGE*
  //(cr_input_valid_realigned_combos): Cover all combinations of realigned versions of the 
  // input valid signals
  
  //*COVERAGE*
  //(cr_valid_realigned_X_embed_combos): Cover all combinations of realigned versions of the 
  // input valid signals
   
  //*COVERAGE*
  //(cp_lreq_w_shifted): Cover the case where there is a link request present
  //from the cs generator but the data is shifted and we are currently out of
  //packet meaning it will need to be selected.

  //*ASSERTION*
  //(ap_dmu_valid_illegal): PTM_valid can never be 2'b01.

  //*COVERAGE*
  //(cr_lreq_X_advance):  Cross all combinations of PTS_lreq with advance 
  //(cr_sop_X_advance):  Cross all combinations of PTS_sop with advance 

  //*COVERAGE*
  //(cr_ccompreq_X_inpkt): See a clock compensation request occur in and out
  //of a packet.

  //*COVERAGE*
  //(cr_ccompreq_X_cs): See a clock compensation request occur when a control
  //symbol needs to be sent.

  //*COVERAGE*
  //(cp_ccomp_w_eop): See a ccomp request occur on an EOP

  //*COVERAGE*
  //(cp_ccomp_w_eop_m1): See a ccomp request occur one cycle before EOP

  //*COVERAGE*
  //(cp_ccomp_w_eop_p1): See a ccomp request occur one cycle after EOP

  //*COVERAGE*
  //(cp_ccomp_w_sop): See a ccomp request occur on SOP
  
  //*COVERAGE*
  //(cp_ccomp_w_sop_m1): See a ccomp request occur one cycle before SOP

  //*COVERAGE*
  //(cp_ccomp_w_sop_p1):  See a ccomp request occur one cycle after SOP

  //*COVERAGE*
  //(cp_ccomp_w_b2b_sop_eop): See a ccomp request occur on EOP followed by an
  //SOP

  //*ASSERTION*
  // (ap_no_ending_cs_on_eop0/ap_no_ending_cs_on_eop1): When an EOP is detected there 
  // must be a control symbol ready to terminate the packet with
  // }}} end Data Mux Control Logic

  // {{{ Register Outputs
  //Dont include a reset on non-control buses
  always @(posedge phy_clk) begin
    if (PTR_ptm_advance) begin
      PTM_data     <= #TCQ data_realigned;
      PTM_charisk  <= #TCQ charisk_realigned;
    end
  end

  wire accepted_lreq = PTS_lreq && PTR_pts_advance;

  //Drive the control which requires a reset
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PTM_tx_early_valid  <= #TCQ 0;
      PTM_tx_early_lreq   <= #TCQ 0;
      PTM_valid           <= #TCQ 0;
      PTM_send_lreq       <= #TCQ 0;
    end else begin
      if (PTR_ptm_advance) begin
        PTM_tx_early_valid  <= #TCQ valid_realigned;
        PTM_tx_early_lreq   <= #TCQ accepted_lreq;
        PTM_valid           <= #TCQ valid_realigned;
        PTM_send_lreq       <= #TCQ accepted_lreq;
      end
    end
  end
  // }}} end Register Outputs

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2010 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/phy/ollm_tx/srio_gen2_v4_1_16_ollm_tx_ready_gen.v#1 $
//----------------------------------------------------------------------
//
// OLLM_TX_READY_GEN
// Description:
// This module generates the advance signal to each stage in the OLLM
//
// Hierarchy:
// PHY_TOP
//    |___OLLM_TX_TOP
//             |_____OLLM_TX_READY_GEN <-- this module
//             |_____OLLM_TX_BUF
//             |_____OLLM_TX_PKT_ASSEMBLY
//             |_____OLLM_TX_CS_GEN
//             |_____OLLM_TX_DATA_MUX
//             |_____OLLM_TX_OPLM  
// ---------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_ollm_tx_ready_gen
  #(
    parameter TCQ         = 100 
  )
  (
    // {{{ Port Declarations
    // System Signals
    input               phy_clk,              // PHY interface clock
    input               phy_rst,              // Reset for PHY clock Domain

    // TX Buffer Interface
    output wire         PTR_phyt_tready,      // Ready to the buffer interface
    
    // OLLM TX Buf Interface
    input               PTB_stall,            // Stall from the OLLMTX BUF module
    output wire         PTR_ptb_advance,      // Advance Indicator to the OLLMTX BUF

    // OLLM TX OPLM Interface
    input               PTP_stall,            // Stall from the OLLMTX OPLM module
    output wire         PTR_ptp_advance,      // Advance Indicator to OLLMTX OPLM

    // OLLM TX Data Mux Interface
    input               PTM_pta_stall,        // Stall from the Data Mux to PA
    input               PTM_pts_stall,        // Stall from the Data Mux to CS Gen
    output wire         PTR_ptm_advance,      // Advance Indicator to the Data Mux

    // OLLM TX Packet Assembly Interface
    input               PTA_in_packet,        // Early in packet indicator
    input               PTA_stall,            // Stall from Packet Assembly 
    output wire         PTR_pta_advance,      // Advance Indicator to the PA

    // OLLM TX Control Symbol Interface
    input               PTS_stall,            // Stall from CS Generator 
    output wire         PTR_pts_advance       // Advance Indicator to the CS Gen
    // }}} end Port Declarations
  );                  
  
  // {{{ Wire Declarations
  reg   phy_rst_q = 1;
  // }}} end wire declarations
  
  // {{{ Register Reset
  // Must register the reset before use
  always @(posedge phy_clk) begin
    phy_rst_q <= #TCQ phy_rst;
  end
  // }}} end Register Reset

  // Advance each module if the modules before it are ready to accept it
  // When a module indicates to stall all stages before that module must also
  // stall. The Buffer has the additional requirement that the link must be
  // initialized before packets can be transmitted. 
  // OLLM TX Stages Order:
  // BUF -> PKT_ASSEMBLY -> DATA_MUX -> OPLM
  //        CS_GEN
  assign PTR_ptm_advance = !PTP_stall;
  assign PTR_pts_advance = !PTP_stall && !PTM_pts_stall;
  assign PTR_pta_advance = !PTP_stall && !(PTS_stall && PTR_pts_advance) && !PTM_pta_stall;
  assign PTR_ptb_advance = !PTP_stall && !PTA_stall && 
                           !(PTS_stall && PTR_pts_advance) && !PTM_pta_stall;
  assign PTR_phyt_tready = !PTP_stall && !PTA_stall && 
                           !PTB_stall && !(PTS_stall && PTR_pts_advance) && !PTM_pta_stall;

  // The stall to the OPLM module is the same as to the data mux
  assign PTR_ptp_advance = PTR_ptm_advance;

  //*COVERAGE*
  // (cr_advance_stages): Cover all the combinations of advance indicators from 
  // each stage of the OLLM TX pipeline.

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2010 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/phy/ollm_tx/srio_gen2_v4_1_16_ollm_tx_buf.v#1 $
//----------------------------------------------------------------------
//
// OLLM_TX_BUF_AXI
// Description:
// This module is the TX Buffer AXI Interface of the OLLM TX design. It 
// is responsible for:
// 1. swizzling the axi formatting to SRIO packet format
// 2. registering incoming data from the TX Buffer
// 3. generating sideband signals to the rest of the design
// 4. generating the packet ID and drive next_fm to the TX Buffer
// 5. generating the CRC value as data is accepted 
//
// Hierarchy:
// PHY_TOP
//    |___OLLM_TX_TOP
//             |_____OLLM_TX_READY_GEN
//             |_____OLLM_TX_BUF  <-- this module
//             |_____OLLM_TX_PKT_ASSEMBLY
//             |_____OLLM_TX_CS_GEN
//             |_____OLLM_TX_DATA_MUX
//             |_____OLLM_TX_OPLM
// ---------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_ollm_tx_buf
  #(
    parameter TCQ         = 100,
    parameter IDLE1       = 1,  // Include the IDLE1 Sequence Logic
    parameter IDLE2       = 0,  // Include the IDLE2 Sequence Logic
    parameter SWITCH_MODE = 0)  // Include Switch Mode Support 
  (
    // {{{ Port Declarations
    // System Signals
    input               phy_clk,              // PHY interface clock
    input               phy_rst,              // Reset for PHY clock Domain
    
    // TX Buffer Interface Signals
    input               BT_phyt_tvalid,       // Valid data indicator
    input               PT_phyt_tready,       // Destination Ready
    input       [63:0]  BT_phyt_tdata,        // Packet for transfer
    input       [7:0]   BT_phyt_tkeep,        // Byte Enable for transferred packet
    input               BT_phyt_tlast,        // Last DW of incoming packet
    input       [7:0]   BT_phyt_tuser,        // {1'b0, SKIP_CRC, 2'h00, VC[1:0], CRF, SRC_DSC}
    output reg  [5:0]   PTB_phy_next_fm,      // The next expected frame's ID
    output reg          PTB_phy_rewind,       // Holds PR_rewind high as long as we 
                                              //  are killing a packet 
    // User Global Interface
    input               UG_phy_link_reset,    // Reset the link via control symbols

    // OLLM TX Packet Assembly Interface
    output reg  [5:0]   PTB_next_fm,          // Next ack ID for packets
    output wire         PTB_sop_d,            // One cycle early version of SOP
    output reg          PTB_sop,              // SOP
    output reg          PTB_eop,              // EOP
    output reg          PTB_src_disc,         // Source Disconnect (for STOMP) // cr 800810, stomp
    output reg          PTB_valid,            // Valid Cycle
    output wire         PTB_valid_d,          // Valid Cycle - unregistered
    output reg  [63:0]  PTB_data,             // Data
    output reg  [3:0]   PTB_keep,             // Strobe
    output reg          PTB_vc,               // VC for this packet
    output reg          PTB_crf,              // CRF for this packet
    output reg          PTB_in_packet,        // Indicates in a packet
    output reg          PTB_skip_final_crc,   // Indicates to skip final CRC insertion
    output reg  [15:0]  PTB_crc64,            // The current CRC value 
    output reg  [15:0]  PTB_crc48,            // The current CRC value 
    output reg  [15:0]  PTB_crc32,            // The current CRC value 
    output reg  [15:0]  PTB_crc16,            // The current CRC value 
    output reg          PTB_insert_mid_crc,   // Insert the mid CRC
    output reg          PTB_mid_crc_inserted, // A mid CRC was inserted

    // OLLM RX Interface
    input               PR_rewind,            // Indicates a rewind is in progress
    input       [5:0]   PR_phy_last_ack,      // Last PA received by the PHY core
    output reg          PTB_sample_next_fm,   // Indicates to the ollm rx to sample the next fm
                                              //  value in a rewind scenario.
    input               PR_link_initialized,  // Indicate if link init is obtained                                          
    // OLLM TX CS Generator Inteface
    input               PTS_lreq_sent,        // A rewind LREQ was sent    
    input               PTS_rfr_sent,         // A rewind RFR was sent
    input               PR_send_lreq,         // A LREQ needs to be sent
    input               PR_send_rfr,          // A RFR needs to be sent
    output reg          PTB_link_reset,       // Send a LREQ/reset-device cs

    // OPLM TX Interface Signals
    input               PP_port_initialized,  // Indicates the port is initialized
    input               PP_idle2_selected,    // Indicates the operating idle mode

    // PHY Config Interface Signals
    input               PC_load_ackids,       // Indication to load Pnext_fm into phy_next_fm
    input       [5:0]   PC_next_fm,           // Value to load into phy_next_fm when

    // OLLM TX Ready Generator Interface
    output reg          PTB_stall,            // Stall from this module
    input               PTR_ptb_advance       // Advance this module
    // }}} end Port Declarations
  );          

  // {{{ Local Parameters
  localparam VC       = 2; // the VC bit of the user bus
  localparam CRF      = 1; // the CRF bit of the user bus
  localparam SRC_DSC  = 0; // the SRC_DSC bit of the user bus
  localparam SKIP_CRC = 6; // the SKIP_CRC bit of the user bus

  // When in IDLE2 mode, ack id's are 6 bits; for IDLE1 mode only 5 bits
  localparam ID_WIDTH = (IDLE2) ? 6 : 5;
  // }}} end Local Parameters

  // {{{ Wire Declarations
  reg           phy_rst_q = 1;

  // Registered inputs from the buffer interface 
  // Stage 1 of this module

  /*
  reg   [5:0]   next_fm_dd;
  reg           ready_dd;          
  reg           valid_dd;          
  reg   [63:0]  data_dd;          
  reg   [7:0]   keep_dd;         
  reg   [7:0]   user_dd;        
  reg           last_dd;       
*/


  wire   [5:0]   next_fm_dd;
  wire           ready_dd;          
  wire           valid_dd;          
  wire   [63:0]  data_dd;          
  wire   [7:0]   keep_dd;         
  wire   [7:0]   user_dd;        
  wire           last_dd;   

  // Registered versions of the phyt_t* signals.
  // Stage 2 of this module before registered outputs
  reg   [5:0]   next_fm_d;
  reg           in_packet_d;          
  reg   [63:0]  data_d;
  reg   [7:0]   last_valid_data_d;
  reg   [3:0]   keep_d;
  reg           sop_d;
  reg           eop_d;
  reg           valid_d;
  reg           src_disc_d; // cr 800810, stomp
  reg           vc_d;
  reg           crf_d;
  reg           skip_final_crc_d;
  reg           max_pkts_stall;     // Stall when no more ack IDs are available
  wire          phyt_active;        // active beat on the PHYT interface
  wire          sop_on_rewind;      // Indicates a SOP on the first rewind beat
  reg           ptb_phy_rewind_q;   // registered PTB_phy_rewind
  wire          phyt_last_active;   // active last beat on the PHYT interface
  wire  [63:0]  swizzled_data_dd;   // SRIO format of data swizzled from AXI format
  wire  [3:0]   swizzled_keep_dd;   // SRIO format of keep swizzled from AXI format 
                                    //  and reduced to 4 bits from 8
  wire          active_cycle_dd;    // indicates valid_dd and phyt_tready are both asserted
  wire          sop_active_dd;      // SOP was detected on the phyt_t* signals
  wire          eop_active_dd;      // EOP was accepted by packet assembly 
  reg           eop_active_d;       // Registered eop_active_dd
  wire          flush_pipe;         // Indicates to flush out this module
  wire          flush_needed;       // A flush needs to occur in this module
  reg           kill_current_pkt;   // Kill the current transmitting pkt
  wire          phyt_active_dd;     // active cycle in stage 1 of this module
  // }}} end Wire Declarations

  // {{{ Register Reset
  // Must register the reset before use
  always @(posedge phy_clk) begin
    phy_rst_q <= #TCQ phy_rst;
  end  
  // }}} end Register Reset

  // {{{ Stage 1 
  // On a rewind scenario, and LREQ or RFR will only be sent
  // at the end of a packet. If anything is leftover in this
  // module it needs to be flushed. specifically small and single
  // cycle packets which will fit in this module completely
  assign flush_pipe = PTS_lreq_sent || PTS_rfr_sent || (!flush_needed && PTB_phy_rewind);

  // In the case of a short rewind we need to hold rewind until the flush
  // occurs
  assign flush_needed = (PR_send_lreq && !PTS_lreq_sent) || 
                        (PR_send_rfr && !PTS_rfr_sent);

  // Register TX Buffer Interface Signals Before Use 
  // This will ease timing between cores.

  // Register Control Buses
  // Dont need a reset on the non-control buses
  
  /*
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      next_fm_dd <= #TCQ 0;
      valid_dd   <= #TCQ 0;
      ready_dd   <= #TCQ 0;
      last_dd    <= #TCQ 0;

    // Clear out the pipe if a new packet is started an a flush needs to occur
    // or when flush_pipe asserts
    end else if (flush_pipe) begin
      next_fm_dd <= #TCQ 0;
      valid_dd   <= #TCQ 0;
      ready_dd   <= #TCQ 0;
      last_dd    <= #TCQ 0;

    end else if (PTR_ptb_advance) begin
      data_dd     <= #TCQ BT_phyt_tdata;
      keep_dd     <= #TCQ BT_phyt_tkeep;
      user_dd     <= #TCQ BT_phyt_tuser; 
      next_fm_dd  <= #TCQ PTB_phy_next_fm;
      valid_dd    <= #TCQ BT_phyt_tvalid;
      ready_dd    <= #TCQ PT_phyt_tready;
      last_dd     <= #TCQ BT_phyt_tlast;
    end
  end  
*/

      assign data_dd     =  BT_phyt_tdata;
      assign keep_dd     =  BT_phyt_tkeep;
      assign user_dd     =  BT_phyt_tuser; 
      assign next_fm_dd  =  PTB_phy_next_fm;
      assign valid_dd    =  BT_phyt_tvalid;
      assign ready_dd    =  PT_phyt_tready;
      assign last_dd     =  BT_phyt_tlast;

  //*ASSERTION*
  //(ap_single_cycle_keep): For a single cycle packet the strobe will 
  //only ever indicate 5 or 7 bytes. 
  // }}} end Stage 1 

  // {{{ Generate Sideband Signals
  //generate active signals based on readys and valids
  assign active_cycle_dd = valid_dd && ready_dd;
  
  // SOF occurs on the first valid cycle after an EOF
  assign sop_active_dd = ((!in_packet_d && valid_dd) || (eop_active_d && valid_dd)) &&
                         active_cycle_dd;

  wire flush_stage_d = (flush_needed && !PTB_in_packet) || flush_pipe;

  // Capture the SKIP_CRC, VC, and CRF bits only on SOF
  // to hold for the duration of this packet. Dont clear on a rewind
  // since it will reset on the next packet anyway
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      vc_d             <= #TCQ 0;
      crf_d            <= #TCQ 0;
      skip_final_crc_d <= #TCQ 0;
    end else begin
      if (flush_stage_d) begin
        vc_d             <= #TCQ 0;
        crf_d            <= #TCQ 0;
        skip_final_crc_d <= #TCQ 0;

      end else if (sop_active_dd && PTR_ptb_advance) begin
        vc_d  <= #TCQ user_dd[VC];
        crf_d <= #TCQ user_dd[CRF];

        // If switch mode is enabled we need to sample the skip crc bit as
        // well; if we are not in switch mode this bit does not exists.
        // When sampling, for single cycle packets we need to check the
        // the strobe as well to validate that bit.
        skip_final_crc_d <= #TCQ (!SWITCH_MODE) ? 0 :
                                  (user_dd[SKIP_CRC] && keep_dd[SKIP_CRC]); 
      end
    end
  end

  //*COVERAGE*
  //(cp_vc_changed_across_dsc):Cover a change in vc across a discontinued packet
  
  //*COVERAGE*
  //(cp_crf_changed_across_dsc):Cover a change in crf across a discontinued packet
  
  //*COVERAGE*
  //(cp_skip_crc_changed_across_dsc):Cover a change in skip_crc across a discontinued packet

  // Generate in_packet
  // In packet lasts from the detection of SOP to EOP the acceptance of the
  // eof beat. Clear this signal on a rewind if we were in packet
  assign eop_active_dd = last_dd && active_cycle_dd;
 
  //Register eop_active_dd to detect a new sop for single cycle packets
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      eop_active_d <= #TCQ 0;
    end else begin
      if (flush_stage_d) begin
        eop_active_d <= #TCQ 0;

      end else if (PTR_ptb_advance) begin
        eop_active_d <= #TCQ eop_active_dd;
      end
    end
  end

  // This signal is used in the data mux to determine dead beats within
  // packets
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      in_packet_d <= #TCQ 0;
    end else begin
      if (flush_stage_d) begin
        in_packet_d <= #TCQ 0;

      end else if (sop_active_dd && PTR_ptb_advance) begin
        in_packet_d <= #TCQ 1;

      end else if (eop_active_d && PTR_ptb_advance) begin
        in_packet_d <= #TCQ 0;
      end
    end
  end
  // }}} end Generate Sideband Signals

  // {{{ Stage 2
  // Swizzle the incoming data and strobe from AXI Streaming Format
  // to SRIO Packet format and register these inputs
  assign swizzled_data_dd = {data_dd[7:0],   data_dd[15:8],  data_dd[23:16], 
                             data_dd[31:24], data_dd[39:32], data_dd[47:40], 
                             data_dd[55:48], data_dd[63:56]};

  // Strip the strobe down to only 4-bits since we know the only valid
  // combinations are:
  // 8'b1000_0000, 8'b1110_0000, 8'b1111_1000, 8'b1111_1110
  assign swizzled_keep_dd = {keep_dd[0], keep_dd[2], keep_dd[4], keep_dd[6]};

  //Register the captured signals 
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      eop_d     <= #TCQ 0;
      valid_d   <= #TCQ 0;
      sop_d     <= #TCQ 0;
      src_disc_d<=  #TCQ 0; // cr 800810, stomp

    end else begin
      if (flush_stage_d) begin
        eop_d     <= #TCQ 0;
        valid_d   <= #TCQ 0;
        sop_d     <= #TCQ 0;
	    src_disc_d<=  #TCQ 0; // cr 800810, stomp 

      // Update this interface whenever it has been accepted into packet assembly
      end else if (PTR_ptb_advance) begin
        data_d    <= #TCQ swizzled_data_dd;
        keep_d    <= #TCQ swizzled_keep_dd;
        eop_d     <= #TCQ active_cycle_dd && last_dd;
	    src_disc_d<= #TCQ user_dd[SRC_DSC]; // cr 800810, stomp
        valid_d   <= #TCQ active_cycle_dd;
        sop_d     <= #TCQ sop_active_dd;
      end
    end
  end

  // Hold the last valid data_d byte for the crc logic
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      last_valid_data_d <= #TCQ 0;
    end else begin
      if (flush_stage_d) begin
        last_valid_data_d <= #TCQ 0;
      end else if (active_cycle_dd && PTR_ptb_advance) begin
        last_valid_data_d <= #TCQ swizzled_data_dd[7:0];
      end
    end
  end


  //Assign the output wire
  assign PTB_sop_d = sop_d;
  // }}} end Stage 2

  // {{{ Stage 3
  // Flush out this stage on a rewind or a valid SOP is going to propigate
  // during a rewind
  wire flush_last_stage = (flush_needed && !PTB_in_packet) || flush_pipe;

  // Dive to Packet Assembly
  // Register the outputs to be in sync with the 2 stage CRC
  // Do not reset data to save resources
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PTB_eop             <= #TCQ 0;
      PTB_valid           <= #TCQ 0;
      PTB_in_packet       <= #TCQ 0;
      PTB_sop             <= #TCQ 0;
      PTB_vc              <= #TCQ 0;
      PTB_crf             <= #TCQ 0;
      PTB_skip_final_crc  <= #TCQ 0;
      PTB_src_disc        <= #TCQ 0; // cr 800810, stomp
    end else begin 
      if (flush_last_stage) begin
        PTB_eop       <= #TCQ 0;
        PTB_valid     <= #TCQ 0;
        PTB_in_packet <= #TCQ 0;
        PTB_sop       <= #TCQ 0;
	PTB_src_disc  <= #TCQ 0;// cr 800810, stomp

      // Update this interface whenever it has been accepted into packet assembly
      end else if (PTR_ptb_advance) begin
        PTB_data            <= #TCQ data_d;
        PTB_keep            <= #TCQ keep_d;
        PTB_eop             <= #TCQ eop_d;
        PTB_src_disc        <= #TCQ src_disc_d && eop_d; // cr 800810, stomp
        PTB_valid           <= #TCQ valid_d;
        PTB_in_packet       <= #TCQ in_packet_d;
        PTB_sop             <= #TCQ sop_d;
        PTB_vc              <= #TCQ vc_d;
        PTB_crf             <= #TCQ crf_d;
        PTB_skip_final_crc  <= #TCQ skip_final_crc_d;
      end
    end
  end
  // This signal is used to improve performance in the packet assembly block.
  // Don't stall back to the buffer if we see a well-placed dead cycle arriving.
  assign PTB_valid_d = valid_d;

  wire active_pipe = phyt_active || (phyt_active_dd && !last_dd) || 
                    (in_packet_d && !phyt_active_dd && !eop_d);

  assign sop_on_rewind = PTB_phy_rewind && !ptb_phy_rewind_q && BT_phyt_tvalid && !PT_phyt_tready;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      kill_current_pkt <= #TCQ 0;

    // On last whatever pkt we were in is complete and stall back to the
    // buffer now.
    end else if (phyt_last_active) begin
      kill_current_pkt <= #TCQ 1'b0;

    // Keep killing the current packet as long as rewind is asserted and we
    // are in packet
    end else if ((active_pipe && PTB_phy_rewind) || sop_on_rewind) begin
      kill_current_pkt <= #TCQ 1'b1;
    end
  end

  //*COVERAGE*
  //(cp_kill_current_pkt_on_last): kill_current_pkt asserts on the last cycle
  //of a packet

  //*COVERAGE*
  //(cp_kill_current_pkt_on_first): kill_current_pkt asserts on the first cycle
  //of a packet

  //*COVERAGE*
  //(cp_kill_current_pkt_on_valid): kill_current_pkt asserts on a valid cycle
  //of a packet which is not the first or the last

  //*COVERAGE*
  //(cp_kill_current_pkt_on_single): kill_current_pkt asserts on a single cycle
  //packet
  // }}} end Stage 3 

  // {{{ Packet ID Generator
  // Generate the next packets ACK ID value and the next_fm 
  // value to report to the TX Buffer
  // IPCV -
  // need to look directly at the non-registered input in order 
  // for the next fm signal to update directly after last.
  assign phyt_active      = BT_phyt_tvalid && PT_phyt_tready;
  assign phyt_last_active = phyt_active && BT_phyt_tlast;
  wire   idle1_rollover   = !PP_idle2_selected && (&PTB_phy_next_fm[4:0]);
  wire   rewind_rollover  = !PP_idle2_selected && (&PR_phy_last_ack[4:0]);

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PTB_phy_next_fm <= #TCQ 0;

    end else begin
      // Reload the id when indicated by the PHY config
      if (PC_load_ackids) begin
        // Do not load a higher value than is allowed for that idle mode
        PTB_phy_next_fm <= #TCQ (!PP_idle2_selected) ? {1'b0,PC_next_fm[4:0]} : PC_next_fm;
      
        // On a rewind load the next id to be last_ack +1
      end else if (PTB_phy_rewind) begin
        if (phyt_last_active && !flush_last_stage) begin
          PTB_phy_next_fm <= #TCQ (idle1_rollover) ? 0 : PTB_phy_next_fm + 1'b1;
        end else if (flush_pipe) begin
          PTB_phy_next_fm <= #TCQ (rewind_rollover) ? 0 : PR_phy_last_ack + 1'b1;
        end

      // Increment the ack id at the end of every packet when that last beat
      // was accepted.
      end else if (phyt_last_active) begin
        PTB_phy_next_fm <= #TCQ (idle1_rollover) ? 0 : PTB_phy_next_fm + 1'b1;
      end
    end
  end

  // When a rewind occurs the OLLM RX needs to know which value was the actual
  // next_fm value. Indicate a sample time which is needed in case the OLLM TX
  // was in packet when rewind asserted.
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PTB_sample_next_fm <= #TCQ 0;
    end else begin
      if (PTB_sample_next_fm) begin
        PTB_sample_next_fm <= #TCQ 0;

      // Only sample at the end of a rewind or after a valid last beat
      end else if (phyt_last_active && !flush_last_stage) begin
        PTB_sample_next_fm <= #TCQ 1;
      end
    end
  end

  //Register the next frame from the phyt interface to stay in sync
  //with the data to packet assembly
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      next_fm_d     <= #TCQ 0;
      PTB_next_fm   <= #TCQ 0;
    end else begin
      if (PTR_ptb_advance) begin
        next_fm_d     <= #TCQ next_fm_dd;
        PTB_next_fm   <= #TCQ next_fm_d;
      end
    end
  end

  //*COVERAGE*
  //(cp_ackid_rollover_idle2): the ack id counter rolls over in idle2 mode

  //*COVERAGE*
  //(cp_ackid_rollover_idle1): the ack id counter rolls over in idle1 mode
  
  // Outstanding Packets Counter
  // The outstanding packets counter maintains the number of PAs 
  // that need to be sent.
  // REQ: req_pt_idle1_32_pkts_outstanding_max
  // REQ: req_pt_idle2_64_pkts_outstanding_max
  reg   [5:0]          last_ack_q;
  reg   [ID_WIDTH-1:0] outstanding_pkts;

  // Only two bits are used because this is only allowed to change by 3
  // there are assertions in place to check that
  wire [1:0] last_ack_difference = PR_phy_last_ack - last_ack_q;
  
  // Save the last ack value to monitor a change
  // Out of a reset last_ack will either be all ones for IDLE2 mode, or 
  // all ones except for the upper bit for IDLE1 mode
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      last_ack_q <= #TCQ (IDLE2) ? 6'h3F : 6'h1F;
    end else begin
      last_ack_q <= #TCQ PR_phy_last_ack;
    end
  end

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      outstanding_pkts <= #TCQ 0;

    end else begin
      // On a rewind or a reload condition, no more packets are outstanding
      if (PTB_phy_rewind || PC_load_ackids) begin
        outstanding_pkts <= #TCQ 0;

      end else if (PP_port_initialized) begin
        // Increment the outstanding pkt count everytime we send a packet
        // to the packet assembly
        if (phyt_last_active && (last_ack_difference == 0)) begin
          outstanding_pkts <= #TCQ outstanding_pkts + 1'b1;

        // If an ack occurs when last ack changes decrement by the number of
        // acks minues the pkt just sent
        end else if (phyt_last_active && (last_ack_difference != 0)) begin
          outstanding_pkts <= #TCQ outstanding_pkts - (last_ack_difference - 1);

        // Decrement the outstanding pkt count everytime last ack updates
        // this can only increment by 1 unless there is a rewind
        end else if ((last_ack_difference != 0) && !phyt_last_active) begin
          outstanding_pkts <= #TCQ outstanding_pkts - last_ack_difference;
        end
      end
    end
  end

  //*COVERAGE*
  //(cp_link_drop_outstanding_pkts): See link initialized drop when there are
  //ackids outstanding

  //*COVERAGE*
  //(cp_outstanding_pkts_maxed_idle1): outstanding_pkts reaches 30 in idle1 (31 is not allowed
  // due to the number of ack id values)

  //*COVERAGE*
  //(cp_outstanding_pkts_maxed_idle2): outstanding_pkts reaches 62 in idle2 (63 is not allowed
  // due to the number of ack id values)

  //*COVERAGE*
  //(cp_last_ack_w_eof): last_ack_difference and eop_active_dd are both true

  //*ASSERTION*
  //(ap_outstanding_pkts_rollover): outstanding pkts does not rollover 

  //*ASSERTION*
  //(ap_outstanding_pkts_rollunder): outstanding pkts does not rollunder
 
  //*ASSERTION*
  //(ap_outstanding_pkts_changed): Outstanding packets can only ever change by
  //+/- 1

  //*COVERAGE*
  //(cp_outstanding_pkts_maxed_single_inc): Cover that the outstanding
  //packets counter is maxed and a single cycle packet is seen on the _dd
  //interface.

  //*COVERAGE*
  //(cp_outstanding_pkts_enum): enumerate the values of outstanding pkts
  
  //*COVERAGE*
  //(cr_outstanding_pkts_X_last_ack_jumps): Cross the values of outstanding pkts with 
  // a change in last ack

  //*COVERAGE*
  //(cr_outstanding_pkts_X_rewinds): See a rewind with all combinations of outstanding packets
 
  //*ASSERTION*
  //(ap_stalls_ready): If PTB_stall is asserted PT_phyt_tready must be 0 on the next cycle

  //*ASSERTION*
  //(ap_last_ack_invalid_incr): PR_phy_last_ack never increments by more than 1 out of a rewind

  //*COVERAGE*
  //(cp_port_init_drops_stage1): Cover that port init with valid, sop, and eop in
  //stage1 

  //*COVERAGE*
  //(cp_port_init_drops_stage2): Cover that port init with valid, sop, and eop in
  //stage2

  //*COVERAGE*
  //(cp_port_init_drops_stage3): Cover that port init with valid, sop, and eop in
  //stage3
  
  // When outstanding packets reaches the max allowed, we need to stall
  // incoming data.  
  // for idle2 it is when there is 63 and for idle1 it is 31. the ollm_rx
  // needs one pkt leeway to know if the buffer is full or empty so 62 and 30 
  // are used
  // REQ: req_pt_only_send_free_ackids
  reg  max_pkts_stall_q;

  wire [5:0] outstanding_pkts_max = (PP_idle2_selected) ? 61 : 29;

  always @* begin
    //If we havnt reached the max count, dont stall
    if (outstanding_pkts < outstanding_pkts_max) begin
      max_pkts_stall = 0;

    //Stall when we recieve the max number of packets on last so the next
    //SOP wont be accepted if they are back to back
    end else if (phyt_last_active) begin
      max_pkts_stall = 1;

    end else begin
      max_pkts_stall = max_pkts_stall_q;
    end
  end

  // Latch the max_pkts_stall signal
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      max_pkts_stall_q <= #TCQ 0;
    end else begin
      max_pkts_stall_q <= #TCQ max_pkts_stall;
    end
  end
  
  //*COVERAGE*
  //(cp_ptb_stalled): PTB_stall crossed with PP_idle2_selected
  // }}} end Packet ID Generator
 
  // {{{ Rewind Generation
  // Propigate the PR_rewind signal to the TX Buffer interface as long as
  // we are killing a packet. If a packet is currently not in progress then
  // this signal will simply be a registered version of PR_rewind signal
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PTB_phy_rewind <= #TCQ 0;

    end else begin
      // Assert when the OLLM RX indicates a rewind condition
      // Extend the pulse of rewind from the ollm rx if we need to have the
      // ollm rx sample the properly value for next_fm (in the case of an in
      // packet rewind). Rewind must remain asserted until the pulse is
      // sampled in order to assure when rewind drops next_fm is last_ack+1
      // (indicated by phyt_last_active && PTB_phy_rewind)
      if (PC_load_ackids || PR_rewind || flush_needed || 
          (kill_current_pkt && !phyt_last_active)) begin
        PTB_phy_rewind <= #TCQ 1'b1;

      // Do not release rewind until any valid data on this interface is cleared.
      end else if ((flush_pipe || !flush_needed) && !PTB_sample_next_fm) begin
        PTB_phy_rewind <= #TCQ 1'b0;
      end
    end
  end

  // register rewind to find the rising edge
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      ptb_phy_rewind_q <= #TCQ 0;
    end else begin
      ptb_phy_rewind_q <= #TCQ PTB_phy_rewind;
    end
  end
  // }}} end Rewind Generation

  // {{{ Stall Generation
  reg rewind_stall;
  reg rewind_stall_q;
  reg link_init_stall;
  reg link_init_stall_q;
  reg link_reset_stall;
  reg link_reset_stall_q;

  // Stall the buffer interface if:
  // 1. we have reached the max number of ack IDs available
  // 2. We are in a rewind and not killing a pkt
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PTB_stall <= #TCQ 1;
    end else begin
      PTB_stall <= #TCQ max_pkts_stall || rewind_stall || link_init_stall || link_reset_stall;
    end
  end

  // On a rewind, if we are in packet, the remainder of the packet is 
  // masked off until last is seen 
  assign phyt_active_dd = ready_dd && valid_dd;

  wire processing_pkt = kill_current_pkt || active_pipe;

  always @* begin
    if ((!PR_rewind && !flush_needed) || sop_on_rewind) begin
      rewind_stall = 1'b0;

    // Dont start a rewind stall if a kill_current_pkt is about to assert
    // or is already asserted
    end else if (!processing_pkt || phyt_last_active) begin
      rewind_stall = 1'b1;

    end else begin
      rewind_stall = rewind_stall_q;
    end
  end  

  // Latch the rewind_stall signal
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      rewind_stall_q <= #TCQ 0;
    end else begin
      rewind_stall_q <= #TCQ rewind_stall;
    end
  end

  // Stall when link init is not asserted only when we are out of packet.
  always @* begin
    if (PR_link_initialized) begin
      link_init_stall = 1'b0;
    end else if (!PR_link_initialized && (phyt_last_active || !active_pipe)) begin
      link_init_stall = 1'b1;
    end else begin
      link_init_stall = link_init_stall_q;
    end
  end
  
  // Latch the rewind_stall signal
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      link_init_stall_q <= #TCQ 0;
    end else begin
      link_init_stall_q <= #TCQ link_init_stall;
    end
  end

  // Sync and Register the UG signal since it is a core input from the user
  reg        phy_link_reset;
  reg [15:0] ug_phy_link_reset_sync;
  reg        ug_phy_link_reset_sync_q;
  reg        ug_phy_link_reset_sync_qq;

  always @(posedge phy_clk or posedge UG_phy_link_reset) begin
    if (UG_phy_link_reset) begin
      ug_phy_link_reset_sync <= #TCQ 16'hFFFF;
    end else begin
      ug_phy_link_reset_sync <= #TCQ {ug_phy_link_reset_sync[14:0], 1'b0};
    end
  end
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      ug_phy_link_reset_sync_q   <= #TCQ 1'b0;
      ug_phy_link_reset_sync_qq  <= #TCQ 1'b0;
      phy_link_reset             <= #TCQ 1'b0;
    end else begin
      ug_phy_link_reset_sync_q   <= #TCQ |ug_phy_link_reset_sync;
      ug_phy_link_reset_sync_qq  <= #TCQ ug_phy_link_reset_sync_q;
      phy_link_reset             <= #TCQ ug_phy_link_reset_sync_qq;
    end
  end
  
  // If UG_phy_link_reset asserts, wait for the current packet to complete 
  // and then stall so LREQ/reset-device control symbols can be sent. We must
  // complete the packet first since the OLLM TX does not kill packets.
  // link_reset control symbols should not be sent until the port is initialized.
  always @* begin
    if (!phy_link_reset) begin
      link_reset_stall = 1'b0;
    end else if (PP_port_initialized && phy_link_reset && (phyt_last_active || !active_pipe)) begin
      link_reset_stall = 1'b1;
    end else begin
      link_reset_stall = link_reset_stall_q;
    end
  end
  
  // Latch the rewind_stall signal
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      link_reset_stall_q <= #TCQ 0;
    end else begin
      link_reset_stall_q <= #TCQ link_reset_stall;
    end
  end

  // Indicate to send a link reset once the pipe is clear and the buffer is
  // stalled.
  wire data_in_pipe = valid_dd || valid_d;
  wire last_out_pipe = PTB_valid && PTR_ptb_advance && PTB_eop;

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PTB_link_reset <= #TCQ 0;
    end else begin
      if (!link_reset_stall_q) begin
        PTB_link_reset <= #TCQ 0;
      end else if ((last_out_pipe || !data_in_pipe) && link_reset_stall_q) begin
         PTB_link_reset <= #TCQ 1;
      end
    end
  end
  
  // }}} end stall generation

  // {{{ CRC Insertion Counter
  // After 10 cycles (80 bytes of data), a MID-CRC needs to be inserted in the data stream
  reg [3:0] mid_crc_ctr;
  reg       insert_mid_crc_d;
  reg       mid_crc_inserted_d;

  // Reset the mid crc ctr logic:
  // 1. on EOP
  // 2. on a link reset
  wire reset_mid_crc_ctr = eop_active_d || flush_stage_d;

  // Insert the mid crc when the ctr reaches 80 bytes of data
  wire assert_insert_mid_crc = (mid_crc_ctr == 9) && !mid_crc_inserted_d && valid_d;
  
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      insert_mid_crc_d   <= #TCQ 0;

    end else begin
      if (PTR_ptb_advance) begin
        if (reset_mid_crc_ctr || (valid_d && insert_mid_crc_d)) begin
          insert_mid_crc_d <= #TCQ 0;
        end else if (assert_insert_mid_crc) begin
          insert_mid_crc_d <= #TCQ 1;
        end
      end
    end
  end

  //*ASSERTION*
  //(ap_insert_mid_crc_inpkt): PTB_insert_mid_crc can only assert in packet

  //*ASSERTION*
  //(ap_inset_mid_crc_flagged): PTB_insert_mid_crc is only asserted when mid_crc_ctr is 9.

  // Set a flag for when the mid crc has been inserted
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      mid_crc_inserted_d   <= #TCQ 0;

    end else if (PTR_ptb_advance) begin
      if (reset_mid_crc_ctr) begin
        mid_crc_inserted_d   <= #TCQ 0;

      // Use a value of 9 so on the correct on the 10th cycle this will be high
      // one cycle for this to register, then one more for the data to register
      // with the crc in it
      end else if (insert_mid_crc_d && valid_d) begin
        mid_crc_inserted_d <= #TCQ 1;
      end
    end
  end

  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      PTB_insert_mid_crc    <= #TCQ 0;
      PTB_mid_crc_inserted  <= #TCQ 0;
    end else begin
      if (PTR_ptb_advance) begin
        PTB_insert_mid_crc    <= #TCQ insert_mid_crc_d;
        PTB_mid_crc_inserted  <= #TCQ mid_crc_inserted_d;
      end
    end
  end
  
  always @(posedge phy_clk) begin
    if (phy_rst_q) begin
      mid_crc_ctr <= #TCQ 0;

    end else if (PTR_ptb_advance) begin
      if (reset_mid_crc_ctr) begin
        mid_crc_ctr <= #TCQ 0;

      end else if (valid_d) begin
        mid_crc_ctr <= #TCQ mid_crc_ctr + 1'b1;
      end
    end
  end

  //*COVERAGE*
  //(cp_crc_rollover): The CRC counter rolls over

  //*COVERAGE*
  //(cp_link_reset_before_crc): A Link Reset occurs before the CRC is inserted

  //*COVERAGE*
  //(cp_link_reset_on_crc): A Link Reset occurs on CRC is insertion

  //*COVERAGE*
  //(cp_link_reset_after_crc): A Link Reset occurs after the CRC is inserted

  //*COVERAGE*
  //(cp_link_reset_sop): A Link Reset occurs on SOP
  
  //*COVERAGE*
  //(cp_link_reset_eop): A Link Reset occurs on EOP

  //*COVERAGE*
  //(cp_link_reset_midpkt): A Link Reset occurs mid-packet
    
  //*COVERAGE*
  //(cp_link_reset_single_cycle): A Link Reset occurs on a single cycle
  // }}} end CRC Insertion Counter

  // {{{ + CRC-16 Generator +
  // Generate the CRC value for the incoming packet. No reset is needed
  // because it resets on every SOF before use.
  reg   [63:0]  crc64_data_d;
  reg   [15:0]  current_crc_d;
  wire  [15:0]  crc16_d;
  wire  [15:0]  crc32_d;
  wire  [15:0]  crc48_d;
  wire  [15:0]  crc64_d;

  always @(posedge phy_clk) begin
    // Reset the CRC to all 1's at the start of every packet
    // on SOP, include the first byte as all 0's for the Ack ID)
    // REQ: req_pt_crc16_init_value
    if (sop_active_dd && PTR_ptb_advance) begin
      crc64_data_d  <= #TCQ {6'b0, user_dd[VC], user_dd[CRF], swizzled_data_dd[63:8]};
      current_crc_d <= #TCQ 16'hFFFF;

    // Following SOP the data will need to be shifted by 1 byte
    // due to the inserted Ack ID
    end else if (active_cycle_dd && PTR_ptb_advance) begin
      current_crc_d <= #TCQ assert_insert_mid_crc || (insert_mid_crc_d && !valid_d) ? 16'b0 : crc64_d;
      crc64_data_d  <= #TCQ {last_valid_data_d, swizzled_data_dd[63:8]};

    end else if (!active_cycle_dd && PTR_ptb_advance && assert_insert_mid_crc) begin
      current_crc_d <= #TCQ 0;
    end
  end

  //*ASSERTION*
  //(ap_crc_all_ones): On the start of a packet the CRC must be all 1's

  // Register the outputs
  // Calculate the value of the CRC for various valid bytes
  // The correct CRC will be choosen during packet assembly
  always @(posedge phy_clk) begin
    if (PTR_ptb_advance) begin
      PTB_crc16 <= #TCQ crc16_d;
      PTB_crc32 <= #TCQ crc32_d;
      PTB_crc48 <= #TCQ crc48_d;
      PTB_crc64 <= #TCQ crc64_d;
    end
  end

  // 16-bit wide Next CRC Combinational Equations
  srio_gen2_v4_1_16_crc16_16 ollm_tx_crc16_16_inst ( 
    .din   (crc64_data_d[63:48]), 
    .cin   (current_crc_d), 
    .crc   (crc16_d) 
  ); 

  // 32-bit wide Next CRC Combinational Equations
  srio_gen2_v4_1_16_crc16_32 ollm_tx_crc16_32_inst ( 
    .din   (crc64_data_d[63:32]), 
    .cin   (current_crc_d), 
    .crc   (crc32_d) 
  ); 

  // 48-bit wide Next CRC Combinational Equations
  srio_gen2_v4_1_16_crc16_48 ollm_tx_crc16_48_inst ( 
    .din   (crc64_data_d[63:16]), 
    .cin   (current_crc_d), 
    .crc   (crc48_d) 
  ); 

  // 64-bit wide Next CRC Combinational Equations
  srio_gen2_v4_1_16_crc16_64 ollm_tx_crc16_64_inst ( 
    .din   (crc64_data_d), 
    .cin   (current_crc_d), 
    .crc   (crc64_d) 
  ); 
  // }}} + end CRC-16 Generator +

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//---------------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/buf/srio_gen2_v4_1_16_buf_top.v#1 $
//---------------------------------------------------------------------------
//
// BUF_TOP
// Description:
// This module instantiates all the submodules of the BUFFER design
//
// Hierarchy:
// BUF_TOP <-- this module
// ---------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)

module srio_gen2_v4_1_16_buf_top
#(
  parameter TCQ         = 100,
  parameter HW_ARCH     = 2,    // {0 - 8} indication of architecture
  parameter REQ_REORDER = 1,    // {0, 1}
  parameter TX_DEPTH    = 32,   // {8, 16, 32}
  parameter RX_DEPTH    = 32,   // {8, 16, 32}
  parameter RX_FC_ONLY  = 0,    // {0, 1}
  parameter UNIFIED_CLK = 0,    // {0, 1}
  parameter MODE_XG     = 5,    // {1, 2, 3, 4, 5, 6}
  parameter WM0         = 3,    // 62 > WM0
  parameter WM1         = 2,    // WM0 > WM1 > WM2
  parameter WM2         = 1,    // WM2 > 0
  parameter IDLE2       = 0,    // IDLE2 sequence support
  parameter EVAL        = 1)    // {0, 1}
(
  // {{{ port declarations
  //SYSTEM Interface
  input             phy_clk,
  input             log_clk,
  input             cfg_clk,
  input             buf_rst,
  input             cfg_rst,

  //LOG TX Interface
  input             LD_buft_tvalid,       //Valid Packet Beat
  output            BT_buft_tready,       //Packet Beat Accepted
  input   [63:0]    LD_buft_tdata,        //Packet Data
  input   [7:0]     LD_buft_tkeep,        //Valid Bytes in this beat, only valid on last
  input             LD_buft_tlast,        //Last Beat
  input   [7:0]     LD_buft_tuser,        //{4'h00, Response, VC, CRF, 1'b0} AXI Compliance Pad
  output            BT_response_only,     //Buffer only has room for Resp Packets

  //PHY TX Interface
  output            BT_phyt_tvalid,       //Valid Data Indicator
  input             PT_phyt_tready,       //Destination Ready
  output  [63:0]    BT_phyt_tdata,        //Packet Data
  output  [7:0]     BT_phyt_tkeep,        //Byte Enable for data, only valid on last
  output            BT_phyt_tlast,        //Last Beat of Packet Data
  output  [7:0]     BT_phyt_tuser,        //{1'b0, SKIP_CRC, 2'b00, VC[1:0], CRF, SRC_DSC}
  output            BT_tx_flow_control,   //TX Flow Control Mode
  input             PC_master_enable,     //Enable Request Transactions
  input             PP_idle2_selected,    //OPLM has trained to use IDLE2 sequence
  input   [5:0]     PR_phy_rcvd_buf_stat, //Buffer Status received from link partner
  input   [5:0]     PR_phy_last_ack,      //Last PA Received by the PHY
  input   [5:0]     PT_phy_next_fm,       //Next Packet's Ack ID
  input             PT_phy_rewind,        //An Errror or Retry Condition

  //LOG RX Interface
  output            BR_bufr_tvalid,       //Valid Packet Beat
  input             LE_bufr_tready,       //Packet Beat Accepted
  output  [63:0]    BR_bufr_tdata,        //Packet Data
  output  [7:0]     BR_bufr_tkeep,        //Valid bytes in this beat, only valid on last
  output            BR_bufr_tlast,        //Last Beat
  output  [7:0]     BR_bufr_tuser,        //{5'h00, VC, CRF, 1'b0}

  //PHY RX Interface
  input             PR_phyr_tvalid,       //Valid Data Indicator
  output            BR_phyr_tready,       //Destination Ready
  input   [63:0]    PR_phyr_tdata,        //Packet Data
  input   [7:0]     PR_phyr_tkeep,        //Byte Enable for Data, only valid on last
  input             PR_phyr_tlast,        //Last DW of Packet Data
  input   [7:0]     PR_phyr_tuser,        //{5'h00, VC, CRF, src_dsc} AXI Compliance Pad
  output  [5:0]     BR_phy_buf_stat,      //Buffer Status from the RX Buffer

  //CONFIGURATION Interface
  input            CF_cfgb_awvalid,       //Write Command Valid
  output           BC_cfgb_awready,       //Write Port Ready
  input   [23:0]   CF_cfgb_awaddr,        //Write Address
  input            CF_cfgb_wvalid,        //Write Data Valid
  output           BC_cfgb_wready,        //Write Port Ready
  input   [31:0]   CF_cfgb_wdata,         //Write Data
  input   [3:0]    CF_cfgb_wstrb,         //Write Data Byte Enables
  output           BC_cfgb_bvalid,        //Write Response Valid
  input            CF_cfgb_bready,        //Write Response Fabric Ready
  input            CF_cfgb_arvalid,       //Read Command Valid
  output           BC_cfgb_arready,       //Read port Ready
  input   [23:0]   CF_cfgb_araddr,        //Read Address
  output           BC_cfgb_rvalid,        //Read Response Valid
  input            CF_cfgb_rready,        //Read response Fabric Ready
  output  [31:0]   BC_cfgb_rdata          //Read Data
  // }}} end ports
);

// added below macro to fix the CR# 735137
// synthesis translate_off 
  // {{{ Catch Bad Parameters
  //Catch any invalid parameter conditions
  initial begin
    //If IDLE2 is not selected then the highest watermark (WM0) can not be
    //higher than 29. This is because the rcvd_buf_stat can only go to 30 in
    //TX Flow Controlso in order to send out packets it needs to be one less
    //than the highest rcvd_buf_stat
    if (!IDLE2 && (WM0 > 29)) begin
      $display("ERROR: Invalid WM0 value selected for the Buffer based on IDLE2=%0d. WM0=%0d",
                IDLE2, WM0);
      $finish;
    end
  end
  // }}}
// synthesis translate_on

  // {{{ wire declarations -----------------
  wire    [5:0]     BC_watermark0;
  wire    [5:0]     BC_watermark1;
  wire    [5:0]     BC_watermark2;
  wire              BC_force_rx_flow;
  wire              buf_log_rst;
  wire              buf_phy_rst;
  // }}} ---------------------------------

   // {{{ Reset Synchronization ------------
    (* ASYNC_REG = "TRUE" *)
   reg [3:0] buf_log_rst_sr;
   always@(posedge log_clk or posedge buf_rst) begin
     if (buf_rst)
       buf_log_rst_sr <= 4'b1111;
     else
       buf_log_rst_sr <= #TCQ {buf_log_rst_sr[2:0], 1'b0};
   end
   assign buf_log_rst = buf_log_rst_sr[3];

    (* ASYNC_REG = "TRUE" *)
   reg [3:0] buf_phy_rst_sr;
   always@(posedge phy_clk or posedge buf_rst) begin
     if (buf_rst)
       buf_phy_rst_sr <= 4'b1111;
     else
       buf_phy_rst_sr <= #TCQ {buf_phy_rst_sr[2:0], 1'b0};
   end
   assign buf_phy_rst = buf_phy_rst_sr[3];
   // }}} ---------------------------------

  srio_gen2_v4_1_16_buf_tx
  #(
    // {{{ Transmit Buffer Instance --------
    .TCQ                  (TCQ),
    .HW_ARCH              (HW_ARCH),
    .RX_FC_ONLY           (RX_FC_ONLY),
    .TX_DEPTH             (TX_DEPTH),
    .REQ_REORDER          (REQ_REORDER),
    .UNIFIED_CLK          (UNIFIED_CLK))
  buf_tx_inst
   (
    .log_clk              (log_clk),
    .phy_clk              (phy_clk),
    .buf_log_rst          (buf_log_rst),
    .buf_phy_rst          (buf_phy_rst),
    .LD_buft_tvalid       (LD_buft_tvalid),
    .BT_buft_tready       (BT_buft_tready),
    .LD_buft_tdata        (LD_buft_tdata),
    .LD_buft_tkeep        (LD_buft_tkeep),
    .LD_buft_tlast        (LD_buft_tlast),
    .LD_buft_tuser        (LD_buft_tuser),
    .BT_response_only     (BT_response_only),

    .BT_phyt_tvalid       (BT_phyt_tvalid),
    .PT_phyt_tready       (PT_phyt_tready),
    .BT_phyt_tdata        (BT_phyt_tdata),
    .BT_phyt_tkeep        (BT_phyt_tkeep),
    .BT_phyt_tlast        (BT_phyt_tlast),
    .BT_phyt_tuser        (BT_phyt_tuser),
    .BT_tx_flow_control   (BT_tx_flow_control),
    .PC_master_enable     (PC_master_enable),
    .PR_phy_rcvd_buf_stat (PR_phy_rcvd_buf_stat),
    .PR_phy_last_ack      (PR_phy_last_ack),
    .PT_phy_next_fm       (PT_phy_next_fm),
    .PT_phy_rewind        (PT_phy_rewind),

    .BC_watermark0        (BC_watermark0),
    .BC_watermark1        (BC_watermark1),
    .BC_watermark2        (BC_watermark2),
    .BC_force_rx_flow     (BC_force_rx_flow)
    // }}} ---------------------------------
   );

  srio_gen2_v4_1_16_buf_rx
  #(
    // {{{ Receive Buffer Instance ---------
    .TCQ                  (TCQ),
    .MODE_XG              (MODE_XG),
    .HW_ARCH              (HW_ARCH),
    .RX_DEPTH             (RX_DEPTH),
    .UNIFIED_CLK          (UNIFIED_CLK),
    .EVAL                 (EVAL))
  buf_rx_inst
   (
    .log_clk              (log_clk),
    .phy_clk              (phy_clk),
    .buf_log_rst          (buf_log_rst),
    .buf_phy_rst          (buf_phy_rst),
    .BR_bufr_tvalid       (BR_bufr_tvalid),
    .LE_bufr_tready       (LE_bufr_tready),
    .BR_bufr_tdata        (BR_bufr_tdata),
    .BR_bufr_tkeep        (BR_bufr_tkeep),
    .BR_bufr_tlast        (BR_bufr_tlast),
    .BR_bufr_tuser        (BR_bufr_tuser),
    .PR_phyr_tvalid       (PR_phyr_tvalid),
    .BR_phyr_tready       (BR_phyr_tready),
    .PR_phyr_tdata        (PR_phyr_tdata),
    .PR_phyr_tkeep        (PR_phyr_tkeep),
    .PR_phyr_tlast        (PR_phyr_tlast),
    .PR_phyr_tuser        (PR_phyr_tuser),
    .BR_phy_buf_stat      (BR_phy_buf_stat)
    // }}} ---------------------------------
   );

  srio_gen2_v4_1_16_buf_cfg_top
  #(
    // {{{ Buffer Config Instance ----------
      .TCQ                (TCQ),
      .TX_DEPTH           (TX_DEPTH),
      .RX_DEPTH           (RX_DEPTH),
      .RX_FC_ONLY         (RX_FC_ONLY),
      .UNIFIED_CLK        (UNIFIED_CLK),
      .WM0                (WM0),
      .WM1                (WM1),
      .WM2                (WM2),
      .IDLE2              (IDLE2))
  buf_cfg_top_inst
   (
      .phy_clk            (phy_clk),
      .buf_phy_rst        (buf_phy_rst),
      .cfg_clk            (cfg_clk),
      .cfg_rst            (cfg_rst),
      .CF_cfgb_awvalid    (CF_cfgb_awvalid),
      .BC_cfgb_awready    (BC_cfgb_awready),
      .CF_cfgb_awaddr     (CF_cfgb_awaddr),
      .CF_cfgb_wvalid     (CF_cfgb_wvalid),
      .BC_cfgb_wready     (BC_cfgb_wready),
      .CF_cfgb_wdata      (CF_cfgb_wdata),
      .CF_cfgb_wstrb      (CF_cfgb_wstrb),
      .BC_cfgb_bvalid     (BC_cfgb_bvalid),
      .CF_cfgb_bready     (CF_cfgb_bready),
      .CF_cfgb_arvalid    (CF_cfgb_arvalid),
      .BC_cfgb_arready    (BC_cfgb_arready),
      .CF_cfgb_araddr     (CF_cfgb_araddr),
      .BC_cfgb_rvalid     (BC_cfgb_rvalid),
      .CF_cfgb_rready     (CF_cfgb_rready),
      .BC_cfgb_rdata      (BC_cfgb_rdata),
      .BT_tx_flow_control (BT_tx_flow_control),
      .BC_watermark0      (BC_watermark0),
      .BC_watermark1      (BC_watermark1),
      .BC_watermark2      (BC_watermark2),
      .PP_idle2_selected  (PP_idle2_selected),
      .BC_force_rx_flow   (BC_force_rx_flow)
    // }}} ---------------------------------
   );

endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/buf/srio_gen2_v4_1_16_buf_tx.v#1 $
//----------------------------------------------------------------------
//
// BUF_TX
// Description:
// This module is the TX path of the BUFFER. It is responsible for the 
// following:
// 1. Receiving Data from the Logical Layer
// 2. Storing and reordering packets until delivery to the Physical Layer
// 3. Clearing acknowledged packets
// 4. Rewinding back to retried packets and retransmitting
//   
// Hierarchy:
// BUF_TOP
//  |______BUF_TX <-- this module
//  |____________BUF_TX_SYNC_UNIT
//  |____________BUF_TX_BRAM_BANK
//  |______BUF_RX
//  |____________BUF_RX_ASYNC_PASSAGE
//  |____________BUF_RX_BRAM_BANK
// ---------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_buf_tx
  #(
    parameter TCQ           = 100,
    parameter HW_ARCH       = 2,           // {0 -8} indication of architecture
    parameter RX_FC_ONLY    = 0,           // {0, 1} When 1, force Receiver Flow Control
    parameter TX_DEPTH      = 32,          // {8, 16, 32}
    parameter REQ_REORDER   = 1,           // {0, 1} When 1, allows requests to be reordered
    parameter UNIFIED_CLK   = 0)           // {0, 1} When 1, use a common clock
   (
    // {{{ port declarations ---------------
    // clocks and resets
    input             log_clk,             // Freerunning Logical Layer clock
    input             phy_clk,             // Freerunning Physical Layer clock
    input             buf_log_rst,         // Synchronous Logical Layer reset
    input             buf_phy_rst,         // Synchronous Physical Layer reset

    // LOG TX Interface
    input             LD_buft_tvalid,       // Valid Packet Beat
    output            BT_buft_tready,       // Packet Beat Accepted
    input      [63:0] LD_buft_tdata,        // Packet Data
    input       [7:0] LD_buft_tkeep,        // Valid Bytes in this beat, only valid on last
    input             LD_buft_tlast,        // Last Beat
    input       [7:0] LD_buft_tuser,        // {3'h0, Response, 1'b0, VC, CRF, 1'b0} AXI Compliance Pad
    output            BT_response_only,     // Buffer only has room for Resp Packets

    // PHY TX Interface
    output reg        BT_phyt_tvalid,       // Valid Data Indicator
    input             PT_phyt_tready,       // Destination Ready
    output reg [63:0] BT_phyt_tdata,        // Packet Data
    output reg  [7:0] BT_phyt_tkeep,        // Byte Enable for data, only valid on last
    output reg        BT_phyt_tlast,        // Last Beat of Packet Data
    output reg  [7:0] BT_phyt_tuser,        // {1'b0, SKIP_CRC, 2'b00, VC, CRF, SRC_DSC} 
    input             PC_master_enable,     // Enable Request Transactions
    input       [5:0] PR_phy_rcvd_buf_stat, // Buffer Status received from link partner
    input       [5:0] PR_phy_last_ack,      // Last PA Received by the PHY
    input       [5:0] PT_phy_next_fm,       // Next Packet's Ack ID
    input             PT_phy_rewind,        // An Errror or Retry Condition
    output reg        BT_tx_flow_control =0,// Indicates TX Flow control

    // Configuration signals
    input       [5:0] BC_watermark0,        // Watermark for Priority 0
    input       [5:0] BC_watermark1,        // Watermark for Priority 1
    input       [5:0] BC_watermark2,        // Watermark for Priority 2
    input             BC_force_rx_flow      // Forces RX Flow control
    // }}} ---------------------------------
   );

  // {{{ local parameters ------------------

  // Tag Length: corresponds to index for packet storage
  localparam       C_TAG_LEN     = TX_DEPTH ==  8 ? 3 :
                                   TX_DEPTH == 16 ? 4 :
                                   TX_DEPTH == 32 ? 5 :
                                   1; // undefined

  // Family string: direct conversion from HW_ARCH, used to instantiate architecture-specific components
  localparam       C_FAMILY    = HW_ARCH == 0 ? "virtex5"  :
                                 HW_ARCH == 1 ? "virtex5"  :
                                 HW_ARCH == 2 ? "virtex6"  :
                                 HW_ARCH == 3 ? "virtex6"  :
                                 HW_ARCH == 4 ? "spartan6"  :
                                 HW_ARCH == 5 ? "artix7"   :
                                 HW_ARCH == 6 ? "kintex7"  :
                                 HW_ARCH == 7 ? "virtex7"  :
                                 HW_ARCH == 8 ? "virtex7"  :
                                 HW_ARCH == 9 ? "zynq"  :
                                 HW_ARCH == 10 ? "ultrascale"  :
                                 HW_ARCH == 11 ? "ultrascale"  :
                                 HW_ARCH == 12 ? "ultrascale"  :
                                 HW_ARCH == 13 ? "ultrascale"  :
                                 HW_ARCH == 14 ? "ultrascale"  :
                                                "undefined";

  localparam       C_TX_FC_TUNER = 0; // used to add additional safety in watermark calc, 0 means no added safety
  localparam [2:0] C_INDEX_LEN   = 6; // smallest power of 2 that can address an entire packet
  localparam [3:0] C_ADDR_LEN    = C_TAG_LEN + C_INDEX_LEN;
  localparam [1:0] RESPONSE_CH   = 2'h0;
  localparam [1:0] REQUEST2_CH   = 2'h1;
  localparam [1:0] REQUEST1_CH   = 2'h2;
  localparam [1:0] REQUEST0_CH   = 2'h3; 

// added below macro to fix the CR# 735137
// synthesis translate_off 
  initial begin
    if (C_TAG_LEN == 1) begin
      $display("ERROR: TX_DEPTH holds an unexpected value in buf_tx");
      $finish;
    end
    if (C_FAMILY == "undefined") begin
      $display("ERROR: HW_ARCH holds an unexpected value in buf_tx");
      $finish;
    end
  end
  // }}} ---------------------------------
// synthesis translate_on

  // {{{ wire declarations -----------------
 
  // synchronized versions of the Logical Layer signals
  // All of these signals are driven by the Synchronization Unit
  // BTS prefix - signifies signals originating from the Transmit Buffer's Sync Unit
  wire [63:0]            bts_tx_data;
  wire                   bts_tx_start;
  wire                   bts_tx_last;
  wire                   bts_tx_valid;
  wire [7:0]             bts_tx_user;
  wire [2:0]             bts_tx_keep;
//  reg                    bt_tx_response = 0;
  wire                   bt_tx_ready;


  // buffer related - all of these signals are used in and around the BRAM Bank
  // BTB prefix - signifies signals originating from the Transmit Buffer's BRAM bank
      // write port
  reg                    bt_bram_we = 0;
  reg  [C_INDEX_LEN-1:0] bram_waddr_l; // lower portion of write address
  reg  [C_TAG_LEN-1:0]   bram_waddr_u; // upper portion of write address
  wire [C_ADDR_LEN-1:0]  bt_bram_waddr = {bram_waddr_u, bram_waddr_l};
  wire                   bram_full;
      // read port
  wire                   bt_bram_rd;
  reg  [C_INDEX_LEN-1:0] bram_raddr_l; // lower portion of read address
  reg  [C_TAG_LEN-1:0]   bram_raddr_u; // upper portion of read address
  wire [C_ADDR_LEN-1:0]  bt_bram_raddr = {bram_raddr_u, bram_raddr_l};
      // read information
  reg  [63:0]            btb_tx_data;
  reg                    btb_tx_start;
  reg                    btb_tx_last;
  reg  [2:0]             btb_tx_keep;
  reg  [1:0]             btb_tx_user;
  wire                   btb_tx_bram_last;


  // acknowledge related - all of these signals are used in and around the
  // ACKID block. All of these signals are specifically used for either rewind
  // events or finally clearing a packet once it gets acknowledged.
  // None of these signals are considered to be part of the main stream.
  reg  [4:0]             local_last_acked;       // internal copy of PR_phy_last_ack, used to clear a packet
  reg  [4:0]             local_next_acked;       // closely matches PT_phy_next_fm, used to rewind to a retried packet
  reg  [4:0]             local_next_acked_delay; // closely matches PT_phy_next_fm, used to rewind to a retried packet
  reg                    load_backup;            // causes the read counters to update
  reg                    load_backup_d;          // D input to above register
  reg                    resp_retry;             // kicks off a priority adjust


  // tag related -
  // All of these signals are used in and around the tag logic, which is used
  // to track locations of packets in memory and recall them when needed.
  reg  [TX_DEPTH-1:0]    master_list;           // overall outstanding list
//  reg  [C_TAG_LEN-1:0]   current_write_tag = 0; // gets next_read_tag
  wire [C_TAG_LEN-1:0]   next_write_tag;        // from free location finder
  reg  [C_TAG_LEN-1:0]   next_read_tag;         // from next packet finder
  reg  [C_TAG_LEN-1:0]   current_ack_tag;       // stored value in ack handler
  wire [C_TAG_LEN-1:0]   current_ack_tag_d;     // D input of above register
    // queue tag outputs - next tag in line to be read for each type of packet
  wire [C_TAG_LEN-1:0]   rs_read_tag;
  wire [C_TAG_LEN-1:0]   r2_read_tag;
  wire [C_TAG_LEN-1:0]   r1_read_tag;
  wire [C_TAG_LEN-1:0]   r0_read_tag;
     // write pointers - these point into the four types of storage queues
  reg  [C_TAG_LEN:0]     wrptr_resp_queue;
  reg  [C_TAG_LEN:0]     wrptr_req2_queue;
  reg  [C_TAG_LEN:0]     wrptr_req1_queue;
  reg  [C_TAG_LEN:0]     wrptr_req0_queue;
     // write enables into storage queues
  wire                   wren_resp_queue;
  wire                   wren_req2_queue;
  wire                   wren_req1_queue;
  wire                   wren_req0_queue;
     // read pointers - these point into the four types of storage queues
  reg  [C_TAG_LEN:0]     rdptr_resp_queue;
  reg  [C_TAG_LEN:0]     rdptr_req2_queue;
  reg  [C_TAG_LEN:0]     rdptr_req1_queue;
  reg  [C_TAG_LEN:0]     rdptr_req0_queue;


  // general-use signals
  wire [3:0]             pending_list;          // masked list of pending queues
  wire [3:0]             raw_pending_list;      // masked list of pending queues
  reg                    buf_phy_rst_q = 1;     // registered physical layer reset
  reg                    buf_phy_rst_qq = 1;    // registered physical layer reset
  reg                    buf_phy_rst_qqq = 1;   // registered physical layer reset
  reg                    buf_log_rst_q = 1;     // registered logical layer reset

  wire                   bt_packet_ack;         // 1 when PHY reports an ACK
  reg                    bt_packet_ack_q;       // 1 when PHY reports an ACK
//  reg  [1:0]             wr_priority;           // priority into queue: queue steering signal
  wire [1:0]             rd_priority;           // priority from queue: for prio adjustment
  reg  [1:0]             rd_queue_select;       // which queue to read from
  reg  [1:0]             rd_queue_select_q;     // registered version of above
  wire [1:0]             backup_queue_update;   // enable for backup counters
  reg                    rd_tag_valid;          // new packet is ready for read
  wire                   rd_tag_ack_d;          // ack back to packet finder
  wire                   rd_tag_ack;            // registered version of above
  reg                    rd_tag_ack_pulse;      // single-cycle pulse of rd_tag_ack_d
  reg                    rd_tag_ack_hold;       // held-over version of rd_tag_ack_d
  wire [4:0]             free_buf_partial_sum;  // used to determine free buffer space in link partner
  reg  [5:0]             link_free_buffer;      // how many packets we can send - based on above signal
  reg                    alt_prio_available;    // mux control for alternative priority
  reg                    alt_prio_available_q;  // mux control for alternative priority
  reg  [C_TAG_LEN-1:0]   tag_marker;            // holds tag of retried packet
  reg  [1:0]             rx_prio_adjust;        // adjusted priority
  reg  [1:0]             tx_prio_adjust = 0;    // adjusted priority
  reg                    transmitting_resp = 0; // 1 when transferring a response
  reg  [1:0]             transmit_enable;       // broad enable signal for a transfer
  reg                    pr_phy_rewind_q;       // registered version of rewind signal
  reg                    bt_phyt_tstart;        // start of packet, made to look like an AXI signal
  wire                   bt_phyt_tlast_d;       // D input of the tlast signal going to phy
  reg  [1:0]             bt_phyt_tvalid_d;      // D input to tvalid signal going to phy
  wire                   bt_phyt_advance;       // indicates when to push or pull the pipeline along

  // }}} ---------------------------------


  // {{{ Reset Structure -----------------

  // by rule, we must register the resets before we use them. This is not a
  // synchronizing circuit but rather a method to reduce fanout on the resets.
  //always @(posedge phy_clk or posedge buf_phy_rst) begin
  always @(posedge phy_clk ) begin
    if (buf_phy_rst) begin
      buf_phy_rst_q   <= #TCQ 1'b1;
      buf_phy_rst_qq  <= #TCQ 1'b1;
      buf_phy_rst_qqq <= #TCQ 1'b1;
    end else begin
      buf_phy_rst_q   <= #TCQ 1'b0;
      buf_phy_rst_qq  <= #TCQ buf_phy_rst_q;
      buf_phy_rst_qqq <= #TCQ buf_phy_rst_qq;
    end
  end
  //always @(posedge log_clk or posedge buf_log_rst) begin
  always @(posedge log_clk ) begin
    if (buf_log_rst)
      buf_log_rst_q <= #TCQ 1'b1;
    else
      buf_log_rst_q <= #TCQ 1'b0;
  end


    // *- ASSERTION (BT_reset_behavior)
    // buf_log_rst and buf_phy_rst must overlap when driven high.

  // }}} ---------------------------------


  // {{{ Synchronization Unit -------
  // This unit ensures safe delivery of data between the clock domains.
  // It also uses a counter to keep track of how many packets are
  // outstanding.
  // BTS - signals originating from the Sync Unit, unless it goes out of the TX buffer.

  srio_gen2_v4_1_16_buf_tx_sync_unit
   #(.TCQ                   (TCQ),
     .C_FAMILY              (C_FAMILY),
     .TX_DEPTH              (TX_DEPTH),
     .UNIFIED_CLK           (UNIFIED_CLK))
   buf_tx_sync_unit_inst
    (.log_clk               (log_clk),
     .phy_clk               (phy_clk),
     .buf_log_rst_q         (buf_log_rst_q),
     .buf_phy_rst_q         (buf_phy_rst_q),

     // LOG clock domain signals
     .LD_buft_tlast         (LD_buft_tlast),
     .LD_buft_tvalid        (LD_buft_tvalid),
     .BTS_buft_tready       (BT_buft_tready),
     .LD_buft_tkeep         (LD_buft_tkeep),
     .LD_buft_tdata         (LD_buft_tdata),
     .LD_buft_tuser         (LD_buft_tuser),
     .BTS_response_only     (BT_response_only), // note intentional name change

     // PHY clock domain signals
     .PC_master_enable      (PC_master_enable),
     .BTS_tx_data           (bts_tx_data),
     .BTS_tx_start          (bts_tx_start),
     .BTS_tx_last           (bts_tx_last),
     .BTS_tx_valid          (bts_tx_valid),
     .BTS_tx_user           (bts_tx_user),
     .BTS_tx_keep           (bts_tx_keep),
     .BT_tx_ready           (bt_tx_ready),
     .BT_packet_ack         (bt_packet_ack)
   );


    // *- COVERAGE (BT_outstanding_packets_enumerate)
    // Internal to buf_tx_sync_unit
    // Enumerate outstanding_packets across all valid values (0 through TX_DEPTH + 16)

    // *- ASSERTION (BT_outstanding_packets_behavior)
    // Internal to buf_tx_sync_unit
    // outstanding packets never increments or decrements by more that 1.

    // *- COVERAGE (BT_outstanding_packets_inc_dec)
    // Internal to buf_tx_sync_unit
    // Show that both the increment and decrement condition happen on the same cycle

    // *- ASSERTION (BT_framing_signals_behavior)
    // There should be one TSTART for every TLAST, one TLAST for every TSTART.

  // }}} end Synchronization Unit ---


  // {{{ Write Port Controller ------

  // buffer write address -
  // We handle the two portions of the address seperately, though they are
  // combined for the buffer.
  // Load the upper portion of the buffer on start-of-packet. It gets the next_write_tag.
  // The lower portion should be cleared by the time the next packet arrives.
  // For that matter, clear the lower portion after end-of-packet. Otherwise, for every
  // write to the buffer, increment the lower portion.
  reg  [C_INDEX_LEN-1:0] bram_waddr_l_q; // registered version of address segment
  reg  [C_TAG_LEN-1:0]   bram_waddr_u_q; // registered version of address segment
  always @(posedge phy_clk) begin
    bram_waddr_l_q <= #TCQ bram_waddr_l;
    bram_waddr_u_q <= #TCQ bram_waddr_u;
  end

  // These are used directly to create the write address.
  always @* begin
    // upper portion (tag) - load a new segment location only on start-of-packet.
    if (bts_tx_start && bt_bram_we)
      bram_waddr_u = next_write_tag;
    else
      bram_waddr_u = bram_waddr_u_q;

    // lower portion (index) clear and increment on start-of-packet
    if (bts_tx_start)
      bram_waddr_l = 0;
    // otherwise, increment beat locations after every valid write enable
    else if (bt_bram_we)
      bram_waddr_l = bram_waddr_l_q + 1;
    else
      bram_waddr_l = bram_waddr_l_q;
  end


  // buffer write enable -
  // when both tready and tvalid signals are asserted, issue a write enable to the buffer.
  always @* begin
    bt_bram_we = bt_tx_ready && bts_tx_valid;
  end


  // destination ready (read enable) -
  // The only time the tx buffer must push back is when there are absolutely
  // no packet locations left in memory. We know when there are no locations
  // when the Free Location Finder indicates so. However, we must also allow
  // the current packet to complete before push-back. So, only examine the
  // full indication outside of a streaming packet.
  reg log_out_of_packet_d;
  reg log_out_of_packet;
  always @* begin
    if (bts_tx_last && bts_tx_valid)
      log_out_of_packet_d = 1'b1;
    else if (!bram_full)
      log_out_of_packet_d = 1'b0;
    else 
      log_out_of_packet_d = log_out_of_packet;
  end
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      log_out_of_packet <= #TCQ 1'b1;
    else
      log_out_of_packet <= #TCQ log_out_of_packet_d;
  end
  // Make sure the read enable remains asserted for at least two cycles
  // after the FIFO is reset by using the qqq of the reset here
  assign bt_tx_ready = !(bram_full && log_out_of_packet || buf_phy_rst_qqq);


    // *- COVERAGE (BT_bram_full_with_small_packets)
    // With back-to-back single-cycle packets, cause the buffer to go full + 1.
    // Duplicate this cover point for a unified and non-unified clock

    // *- ASSERTION (BT_bt_bram_we_behavior)
    // The number of write enables to the block ram should match the number of
    // reads out of the synchronization unit

    // *- ASSERTION (BT_sync_unit_read_enable)
    // Show that the read enable to the synchronization unit will remain
    // asserted even when the BRAM indicates it is full in order to finish a packet.

    // *- ASSERTION (BT_sync_unit_read_enable_assert)
    // The read enable to the synchronization unit will not assert for a new packet
    // if the BRAM is full.

    // *- COVERAGE (BT_back_to_back_into_bram)
    // Cover that the write enable is capable of asserting one cycle after a 
    // TLAST, demonstrating zero-cycle turnaround between packets.

    // *- COVERAGE (BT_bram_waddr_non_zero_reset)
    // Observe a reset when both the upper and the lower portions of the write address are non-zero

  // }}} end Write Port Controller --


  // {{{ Write Pointer Maintenance --

  /*
  // Master List update logic -
  // store the current write tag in order to push into one of the queues.
  // Capture on the first cycle so that next_write_tag can update without interfering.
  always @(posedge phy_clk) begin
    if (bts_tx_start && bt_bram_we)
      current_write_tag <= #TCQ bram_waddr_u;
  end


  // packet type determination -
  // grab the priority of the incoming packet in order to select the proper queue to store into.
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      wr_priority <= #TCQ 2'h0;
    else if (bts_tx_start && bt_bram_we)
      wr_priority <= #TCQ bts_tx_data[7:6];
  end


  // Address Tag storage -
  // write pointer queue maintenance. Issue a write enable on every TLAST
  // assertion. Select the appropriate queue based on priority and type.
  reg eof_event; // single-cycle pulse, one cycle after tlast is written into the buffer.
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      eof_event         <= #TCQ 1'b0;
    else
      eof_event         <= #TCQ bts_tx_last && bt_bram_we;
  end
  always @(posedge phy_clk) begin
    if (bts_tx_start && bt_bram_we)
      bt_tx_response    <= #TCQ bts_tx_user[4];
  end

  */


 wire  [C_TAG_LEN-1:0]   current_write_tag; // gets next_read_tag
 wire [1:0] wr_priority;
 wire eof_event;
 wire bt_tx_response;

  reg [1:0] wr_priority_d; 
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      wr_priority_d         <= #TCQ 2'b0;
    else
      wr_priority_d         <= #TCQ wr_priority;
  end
  reg bt_tx_response_d; 
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      bt_tx_response_d         <= #TCQ 1'b0;
    else
      bt_tx_response_d         <= #TCQ bt_tx_response;
  end

 reg  [C_TAG_LEN-1:0]   current_write_tag_d; // gets next_read_tag
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      current_write_tag_d         <= #TCQ 'b0;
    else
      current_write_tag_d         <= #TCQ current_write_tag;
  end

assign wr_priority =  (bts_tx_start && bt_bram_we) ? bts_tx_data[7:6] : wr_priority_d;
assign eof_event =  bts_tx_last && bt_bram_we; 
assign bt_tx_response = (bts_tx_start && bt_bram_we) ?  bts_tx_user[4] : bt_tx_response_d;
assign current_write_tag = (bts_tx_start && bt_bram_we) ?  bram_waddr_u : current_write_tag_d;


  generate if (REQ_REORDER) begin: four_queue_wren_gen
    assign wren_resp_queue =  bt_tx_response && eof_event;
    assign wren_req0_queue = !bt_tx_response && eof_event && (wr_priority == 0);
    assign wren_req1_queue = !bt_tx_response && eof_event && (wr_priority == 1);
    assign wren_req2_queue = !bt_tx_response && eof_event && (wr_priority[1] == 1); // prio = 2 or 3
  end else                  begin: two_queue_wren_gen
    assign wren_resp_queue =  bt_tx_response && eof_event;
    assign wren_req2_queue = !bt_tx_response && eof_event;
  end
  endgenerate

  // Increment the pointers for every TLAST. Store the current_write_tag, not
  // next_write_tag, as it has already incremented to the next location. When
  // the packet is a response, we must also store the priority for potential bumping.
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      wrptr_resp_queue <= #TCQ 0;
      wrptr_req2_queue <= #TCQ 0;
    end else begin
      if (wren_resp_queue)
        wrptr_resp_queue <= #TCQ wrptr_resp_queue + 1;
      if (wren_req2_queue)
        wrptr_req2_queue <= #TCQ wrptr_req2_queue + 1;
    end
  end

  generate if (REQ_REORDER) begin: four_queue_wrpt_gen
    always @(posedge phy_clk) begin
      if (buf_phy_rst_q) begin
        wrptr_req0_queue <= #TCQ 0;
        wrptr_req1_queue <= #TCQ 0;
      end else begin
      if (wren_req1_queue)
        wrptr_req1_queue <= #TCQ wrptr_req1_queue + 1;
      if (wren_req0_queue)
        wrptr_req0_queue <= #TCQ wrptr_req0_queue + 1;
      end
    end
  end
  endgenerate


    // *- COVERAGE (BT_back_to_back_sequence)
    // Write a series of 3 back-to-back single-cycle packets into BRAM
    // to ensure the master list and Write Pointer logic can keep up.

    // *- COVERAGE (BT_back_to_back_sequence_gap1)
    // Write a series of 3 back-to-back single-cycle packets into BRAM
    // with a gap of one cycle between each one.

    // *- COVERAGE (BT_back_to_back_sequence_gap2)
    // Write a series of 3 back-to-back single-cycle packets into BRAM
    // with a gap of two cycles between each one.

    // *- COVERAGE (BT_priority_3_request)
    // Observe a priority 3 request.

    // *- COVERAGE (BT_current_write_tag_enumerate)
    // Enumerate current_write_tag.

    // *- COVERAGE (BT_wr_priority_cross_packet_type)
    // Cross wr_priority with packet type (response/request).

    // *- COVERAGE (BT_wrptr_resp_queue_enumerate)
    // Enumerate wrptr_resp_queue.

    // *- COVERAGE (BT_wrptr_req0_queue_enumerate)
    // Enumerate wrptr_req0_queue.

    // *- COVERAGE (BT_wrptr_req1_queue_enumerate)
    // Enumerate wrptr_req1_queue.

    // *- COVERAGE (BT_wrptr_req2_queue_enumerate)
    // Enumerate wrptr_req2_queue.

    // *- COVERAGE (BT_wrptr_resp_queue_rollover)
    // Observe that wrptr_resp_queue rolls over

    // *- COVERAGE (BT_wrptr_req0_queue_rollover)
    // Observe that wrptr_req0_queue rolls over

    // *- COVERAGE (BT_wrptr_req1_queue_rollover)
    // Observe that wrptr_req1_queue rolls over

    // *- COVERAGE (BT_wrptr_req2_queue_rollover)
    // Observe that wrptr_req2_queue rolls over

    // *- ASSERT (BT_wren_onehot)
    // only one wren_*_queue signal may be asserted at a time.

  // }}} end Write Pointer Maintenance --


  // {{{ Free Location Finder -------

  // this function is used to find a zero in an 8-bit sequence. It returns
  // a 3-bit value which correlates to the address of the location of the zero.
  function [2:0] quadrant_address_lookup(input [7:0] master_list_quadrant);
  begin
    quadrant_address_lookup[2] = &master_list_quadrant[3:0];
    quadrant_address_lookup[1] = &master_list_quadrant[1:0] &&
                                 (&master_list_quadrant[5:4] || !(&master_list_quadrant[3:2]));
    quadrant_address_lookup[0] = (master_list_quadrant[1:0] == 2'h1)  ||
                                 (master_list_quadrant[3:0] == 4'h7)  ||
                                 (master_list_quadrant[5:0] == 6'h1F) ||
                                 (master_list_quadrant[7:0] == 8'h7F);
  end
  endfunction


  reg  [2:0] address_taga = 0; // 3-bit address pointing to a free location within a quadrant of master_list
  reg  [2:0] address_tagb = 0; // 3-bit address pointing to a free location within a quadrant of master_list
  reg  [2:0] address_tagc = 0; // 3-bit address pointing to a free location within a quadrant of master_list
  reg  [2:0] address_tagd = 0; // 3-bit address pointing to a free location within a quadrant of master_list
  reg        sel_a        = 0; // mux select to pick a quadrant
  reg        sel_b        = 0; // mux select to pick a quadrant
  reg        sel_c        = 0; // mux select to pick a quadrant

  // address tag A finds the first free location (zero) in bits [7:0] of the
  // master list. This creates the lower three bits of the address.
  // In all of the following code, the logic operates as follows:
  // tag[2] - this is the uppermost portion of the 3-bit address. It provides
  // the most coarse information. It determines if the first hole (0) is in
  // the upper or lower half of the 8-bit sequence.
  // tag[1] - If tag[2] differentiates between the upper 4 bits and the lower
  // 4 bits, tag[1] differentiates between two-bit sequences.
  // tag[0] - This determines if the first hole is at an even location:
  // 0, 2, 4, or 6. Combining tag[2:0] gives you a complete address for an
  // 8-bit sequence.
  always @* begin
    address_taga = quadrant_address_lookup(master_list[7:0]);
  end

  // address tag B finds the first free location (zero) in bits [15:8] of the
  // master list. This conditionally creates the lower three bits of the
  // address. If the master list is only 8 bits, this logic will not be
  // created. Instead, this register will hold the initial value of zero,
  // eventually getting optimized away in synthesis.
  // Note the logic is the same as the taga logic, only shifted by +8.
  generate if ((TX_DEPTH == 16) || (TX_DEPTH == 32)) begin: tagb_gen
    always @* begin
      address_tagb = quadrant_address_lookup(master_list[15:8]);
    end

    // generate the upper address bits only if needed. Otherwise, they remain
    // initialized to zero. Generate sel_a when the depth is 16 or 32. In
    // other words, when the depth is 8, there is no need to differentiate
    // between the partial addresses; when sel_a is 0, the first quadrant
    // will be used.
    always @* begin
      sel_a = &master_list[7:0];
    end

  end
  endgenerate

  // address tag C and D finds the first free location (zero) in bits [23:16]
  // and [31:24] respectively of the master list. This conditionally creates
  // the lower three bits of the address. If the master list is only 8 or 16
  // bits, this logic will not be created. Instead, this register will hold
  // the initial value of zero, eventually getting optimized away in synthesis.
  // Note the logic is the same as the taga logic, only shifted by +16 and +24.
  generate if (TX_DEPTH == 32) begin: tagcd_gen
    always @* begin
      address_tagc = quadrant_address_lookup(master_list[23:16]);
      address_tagd = quadrant_address_lookup(master_list[31:24]);
    end

    // generate the upper address bits only if needed. Otherwise, they remain
    // initialized about zero. Generate sel_b and sel_c when the depth is 32.
    always @* begin
      sel_b = &master_list[15:8];
      sel_c = &master_list[23:16];
    end

  end
  endgenerate


  // write address tag -
  // This signal is distributed throughout the write side of the tx buffer 
  // logic. When the length of the write tag is shorter than the assignment,
  // the upper bits will be trimmed off.
  // NOTE- for single-cycle packets to pass without adding delay, we can't
  // register this. This is a critical path.
  assign next_write_tag = !sel_a ? {2'b00, address_taga} :
                          !sel_b ? {2'b01, address_tagb} :
                          !sel_c ? {2'b10, address_tagc} :
                                   {2'b11, address_tagd};


  // Buffer full indication -
  // Because of the optimization of the above logic, there is no indication
  // when the buffer is full. This signal looks broadly if there are no zeros
  // in the master list. This is used to create the destination ready signal
  // to the sync unit.
  assign bram_full = &master_list;

  // }}} end Free Location Finder ---


  // {{{ Master List ----------------

  // The Master List is used to keep track of available packet segments in the
  // buffer memory. When a packet segment is occupied, there will be a 1 in that
  // location. When it finally gets ACKed, that location will be cleared to
  // 0. There will be no status change when the packet is merely sent because
  // the packet may eventually be retried.
  wire [TX_DEPTH-1:0] set_cond; // when asserted, set a bit in master_list
  wire [TX_DEPTH-1:0] clr_cond; // when asserted, clear a bit in master_list
  genvar ml_gen;
  generate for
      (ml_gen = 0; ml_gen < TX_DEPTH; ml_gen = ml_gen + 1) begin: mlist_gen

    // Each bit of the master list is set and cleared independently.
    // Thus, the generate loop.

    // clear on an acknowledge event from the ACK ID Maintenance logic.
    assign clr_cond[ml_gen] = (bt_packet_ack_q && (current_ack_tag_d == ml_gen));

    // set on the TSTART from the Logical Layer/Sync Unit.
    assign set_cond[ml_gen] = bts_tx_start && bt_bram_we && (next_write_tag == ml_gen);

    always @(posedge phy_clk) begin
      if (buf_phy_rst_q)
        master_list[ml_gen] <= #TCQ 1'b0;
      else if (clr_cond[ml_gen])
        master_list[ml_gen] <= #TCQ 1'b0;
      else if (set_cond[ml_gen])
        master_list[ml_gen] <= #TCQ 1'b1;
    end

  end
  endgenerate

    // *- COVERAGE (BT_master_list_set_clear_on_diff_bits)
    // Observe a set and clear on different bits within the master_list

    // *- COVERAGE (BT_master_list_consecutive_clears)
    // Observe back-to-back clears on different bits.

    // *- ASSERTION (BT_master_list_double_set)
    // It is not possible for an already-set bit to be set again without first being cleared.

    // *- ASSERTION (BT_master_list_double_clear)
    // It is not possible for an already-cleared bit to be cleared again without first being set.

    // *- ASSERTION (BT_master_list_set_clear_on_same_bits)
    // It is not possible for a bit to be set and cleared on the same cycle.

    // *- COVERAGE (BT_master_list_full)
    // Observe all bits in master_list are set

    // *- COVERAGE (BT_master_list_goes_empty)
    // Observe all bits are cleared (empty) after all bits are set (full)

    // *- COVERAGE (BT_master_list_one_cold)
    // Observe only one single free spot (zero) in each location of master_list

    // *- COVERAGE (BT_master_list_one_hot)
    // Observe only one single occupied spot (one) in each location of master_list

    // *- COVERAGE (BT_master_list_quadrants_full)
    // Observe each quadrant is full while all others are not

    // *- COVERAGE (BT_master_list_reset)
    // Observe a reset when the master list is not empty

  // }}} end Master List ------------


  // {{{ BRAM Bank ------------------

  // intermediate signals, prior to registering
  // BTB - signals originating from the BRAM bank, unless it goes out of the TX buffer.

  reg [C_ADDR_LEN-1:0]  bt_bram_waddr_q;
  reg                   bt_bram_we_q;
  reg [63:0]            bts_tx_data_q;
  reg  [2:1]            bts_tx_user_q; // odd width labelling for consistency of assignment
  reg                   bts_tx_start_q;
  reg                   bts_tx_last_q;
  reg  [2:0]            bts_tx_keep_q;
  always @(posedge phy_clk) begin
    bt_bram_waddr_q  <= #TCQ bt_bram_waddr;
    bts_tx_data_q    <= #TCQ bts_tx_data;
    bts_tx_user_q    <= #TCQ bts_tx_user[2:1];
    bts_tx_start_q   <= #TCQ bts_tx_start;
    bts_tx_last_q    <= #TCQ bts_tx_last;
    bts_tx_keep_q    <= #TCQ bts_tx_keep;
  end
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      bt_bram_we_q     <= #TCQ 1'b0;
    end else begin
      bt_bram_we_q     <= #TCQ bt_bram_we;
    end
  end

  wire [63:0] btb_tx_bram_data;  // intermediate signals between BRAM and registers
  wire  [1:0] btb_tx_bram_user;  // intermediate signals between BRAM and registers
  wire        btb_tx_bram_start; // intermediate signals between BRAM and registers
  wire  [2:0] btb_tx_bram_keep;  // intermediate signals between BRAM and registers

  srio_gen2_v4_1_16_buf_tx_bram_bank
   #(.TCQ                  (TCQ),
     .C_FAMILY             (C_FAMILY),
     .C_INDEX_LEN          (C_INDEX_LEN),
     .C_ADDR_LEN           (C_ADDR_LEN))
   buf_tx_bram_bank_inst
    (.phy_clk              (phy_clk),
     .buf_phy_rst_q        (buf_phy_rst_q),
     // in from tx buffer
     .BT_bram_waddr        (bt_bram_waddr_q),
     .BT_bram_rd           (bt_bram_rd),
     .BT_bram_raddr        (bt_bram_raddr),
     .BT_bram_we           (bt_bram_we_q),
     // in from synchronization unit
     .BTS_tx_data          (bts_tx_data_q),
     .BTS_tx_user          (bts_tx_user_q),
     .BTS_tx_start         (bts_tx_start_q),
     .BTS_tx_last          (bts_tx_last_q),
     .BTS_tx_keep          (bts_tx_keep_q),
     // out to Physical layer
     .BTB_tx_bram_data     (btb_tx_bram_data),
     .BTB_tx_bram_user     (btb_tx_bram_user),
     .BTB_tx_bram_start    (btb_tx_bram_start),
     .BTB_tx_bram_last     (btb_tx_bram_last),
     .BTB_tx_bram_keep     (btb_tx_bram_keep)
    );

  // use fabric registers instead of BRAM registers.
  // This is a trade-off for performance. We can steal tlast information early
  // this way and still register all the other signals at the BRAM to improve timing.
  // The alternative of using BRAM registers is that there would be two dead cycles
  // between packets instead of one.
// INFO - CFR - we can improve resource count by adding registers to the BRAM
// other than the one that outputs TLAST and removing those fabric registers.
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
     btb_tx_data  <= #TCQ 64'h0;
     btb_tx_user  <= #TCQ 2'h0;
     btb_tx_start <= #TCQ 1'b0;
     btb_tx_last  <= #TCQ 1'b0;
     btb_tx_keep  <= #TCQ 3'h0;
    end else if (bt_phyt_advance) begin
     btb_tx_data  <= #TCQ btb_tx_bram_data;
     btb_tx_user  <= #TCQ btb_tx_bram_user;
     btb_tx_start <= #TCQ btb_tx_bram_start && bt_phyt_tvalid_d[0];
     btb_tx_last  <= #TCQ btb_tx_bram_last && bt_phyt_tvalid_d[0];
     btb_tx_keep  <= #TCQ btb_tx_bram_keep;
    end
  end


    // *- COVERAGE (BT_write_on_tlast)
    // When the memory transitions to full, it is possible to stall the final write into the
    // BRAM. Observe bram_we low when tlast is asserted

  // }}} end BRAM Bank --------------


  // {{{ Response/Request Tags ------

  // declare the memories implicitly. Split the response queue into two
  // memories based on function.
  (* ram_style = "distributed" *) reg  [C_TAG_LEN-1:0]  resp_queue      [0:TX_DEPTH-1];
  (* ram_style = "distributed" *) reg  [1:0]            resp_queue_prio [0:TX_DEPTH-1];
  (* ram_style = "distributed" *) reg  [C_TAG_LEN-1:0]  req2_queue      [0:TX_DEPTH-1];
    // these two get removed when REQ_REORDER = 0
  (* ram_style = "distributed" *) reg  [C_TAG_LEN-1:0]  req1_queue      [0:TX_DEPTH-1];
  (* ram_style = "distributed" *) reg  [C_TAG_LEN-1:0]  req0_queue      [0:TX_DEPTH-1];


  // write-side operation-
  // keep this clean to ensure the we get the structure we actually want (dist ram).
  wire [C_TAG_LEN-1:0]   wrptr_resp_queue_rip = wrptr_resp_queue[C_TAG_LEN-1:0];
  wire [C_TAG_LEN-1:0]   wrptr_req2_queue_rip = wrptr_req2_queue[C_TAG_LEN-1:0];
  always @(posedge phy_clk) begin
    if (wren_resp_queue) begin
      resp_queue[wrptr_resp_queue_rip]      <= #TCQ current_write_tag;
      resp_queue_prio[wrptr_resp_queue_rip] <= #TCQ wr_priority;
    end
  end

  always @(posedge phy_clk) begin
    if (wren_req2_queue)
      req2_queue[wrptr_req2_queue_rip] <= #TCQ current_write_tag;
  end

  generate if (REQ_REORDER) begin: four_queue_write_gen
    wire [C_TAG_LEN-1:0]   wrptr_req0_queue_rip = wrptr_req0_queue[C_TAG_LEN-1:0];
    wire [C_TAG_LEN-1:0]   wrptr_req1_queue_rip = wrptr_req1_queue[C_TAG_LEN-1:0];
    always @(posedge phy_clk) begin
      if (wren_req1_queue)
        req1_queue[wrptr_req1_queue_rip] <= #TCQ current_write_tag;
    end

    always @(posedge phy_clk) begin
      if (wren_req0_queue)
        req0_queue[wrptr_req0_queue_rip] <= #TCQ current_write_tag;
    end
  end
  endgenerate


  // read-side operation-
  // keep this clean to ensure the we get the structure we actually want (dist ram).
  // These four tags will be muxed to create the next read tag.
  wire [C_TAG_LEN-1:0]   rdptr_resp_queue_rip = rdptr_resp_queue[C_TAG_LEN-1:0];
  wire [C_TAG_LEN-1:0]   rdptr_req2_queue_rip = rdptr_req2_queue[C_TAG_LEN-1:0];
  assign rs_read_tag = resp_queue[rdptr_resp_queue_rip];
  assign r2_read_tag = req2_queue[rdptr_req2_queue_rip];

  generate if (REQ_REORDER) begin: four_queue_read_gen
    wire [C_TAG_LEN-1:0]   rdptr_req1_queue_rip = rdptr_req1_queue[C_TAG_LEN-1:0];
    wire [C_TAG_LEN-1:0]   rdptr_req0_queue_rip = rdptr_req0_queue[C_TAG_LEN-1:0];
    assign r1_read_tag = req1_queue[rdptr_req1_queue_rip];
    assign r0_read_tag = req0_queue[rdptr_req0_queue_rip];
  end
  endgenerate

  // priority acquisition
  assign rd_priority = resp_queue_prio[rdptr_resp_queue_rip];


    // *- ASSERTION (BT_resp_queue_prio)
    // wr_priority will never be 0 when wren_resp_queue is asserted

  // }}} end Response/Request Tags --


  // {{{ Priority Adjust ------------
  // Priority adjusting happens when a rewind occurs on a response.
  // Priority bumping due to watermarks is handled elsewhere.

  reg                    tag_search; // set when logic should be searching for a tag
  reg                    tag_set;    // single-cycle pulse, indicates beginning of rewind

  // This logic is used to set the search mechanism.
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      tag_set <= #TCQ 1'b0;
    else
      tag_set <= #TCQ load_backup;
  end

  // enable the searching mechanism. Whenever a rewind occurs, this register
  // will get set, not clearing until we find the packet that we're looking
  // for. This logic enables the priority capturing mechanism.
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      tag_search <= #TCQ 1'b0;
    // enable the searching mechanism one cycle after we have loaded the new
    // counters.
    else if (tag_set && resp_retry)
      tag_search <= #TCQ 1'b1;
    // only clear when we see the appropriate tag arrive from the response
    // queue. The same cycle, another piece of logic will capture the new priority.
    else if ((tag_marker == rs_read_tag) || (bt_phyt_tstart && PT_phyt_tready))
      tag_search <= #TCQ 1'b0;
  end

  // the tag from the ACK logic specifies which one has been retried.
  // NOTE - in this instance, current_ack_tag uses tnext_ack address
  always @(posedge phy_clk) begin
    if (tag_set && resp_retry)
      tag_marker <= #TCQ current_ack_tag;
  end


  // RX flow control priority adjust-
  // Only used in RX flow control. Capture and increment the stored tag.
  // Only increment if the number is less than 3. Also, if the packet has
  // been retried more than once, increment the locally stored value instead
  // of the one coming from the Response Queue.
  // Mux beforehand to ensure we don't create two seperate adders.
  // if alt_prio_available, that means this is not the first time we've rewound on this ackid
  wire [1:0] rx_prio_adjust_input = alt_prio_available ? rx_prio_adjust : rd_priority;
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      rx_prio_adjust <= #TCQ 2'b0;
    end else if (tag_search && (tag_marker == rs_read_tag)) begin
      if (rx_prio_adjust_input < 2'h3) begin
        rx_prio_adjust <= #TCQ rx_prio_adjust_input + 1;
      end else begin
        rx_prio_adjust <= #TCQ rx_prio_adjust_input;
      end
    end
  end


  // Set an indication to tell the Control Signal Drivers to swap in the
  // modified priority.
  always @(posedge phy_clk) begin
    // make sure to only swap in the retried priority but still hold on to the
    // value in case it gets retried a second time.
    if (buf_phy_rst_q)
      alt_prio_available <= #TCQ 1'b0;
    else if (tag_search && &transmit_enable && (tag_marker == rs_read_tag))
      alt_prio_available <= #TCQ 1'b1;
    // NOTE - in this instance, current_ack_tag uses tlast_ack address
    else if (bt_packet_ack_q && (current_ack_tag_d == tag_marker))
      alt_prio_available <= #TCQ 1'b0;
  end
  always @(posedge phy_clk) begin
    alt_prio_available_q <= #TCQ alt_prio_available;
  end


    // *- COVERAGE (BT_bump_priority_again)
    // See the same response packet get retried a second time.
    // tag_search && (tag_marker == rs_read_tag) && alt_prio_available

    // *- COVERAGE (BT_retry_prio_3_response)
    // Issue a retry on a priority 3 response. It should not bump priority.

    // *- COVERAGE (BT_retry_response)
    // Issue a retry on a response other than priority 3.

    // *- COVERAGE (BT_retry_request)
    // Issue a retry on a request packet.

    // *- COVERAGE (BT_original_cross_modified_priority)
    // Observe all legal combinations of original priority and modified priority

  // }}} end Priority Adjust --------


  // {{{ Read Pointer Maintenance ---

  // dedicate registers for the backup of the read pointers
  reg  [C_TAG_LEN:0]    rdptr_backup_resp_queue; // backup counters for rewind event
  reg  [C_TAG_LEN:0]    rdptr_backup_req2_queue; // backup counters for rewind event
    // These two are removed when REQ_REORDER = 0
  reg  [C_TAG_LEN:0]    rdptr_backup_req0_queue; // backup counters for rewind event
  reg  [C_TAG_LEN:0]    rdptr_backup_req1_queue; // backup counters for rewind event

  // Increment the pointers when indicated by the Next Packet Finder. When
  // requested, load the backup values from the alternate counters.
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      rdptr_resp_queue <= #TCQ 0;
      rdptr_req2_queue <= #TCQ 0;
    end else if (load_backup) begin // backup indication - load backup values
        rdptr_resp_queue <= #TCQ rdptr_backup_resp_queue;
        rdptr_req2_queue <= #TCQ rdptr_backup_req2_queue;
    end else if (rd_tag_ack) begin
      if (rd_queue_select_q == RESPONSE_CH)
        rdptr_resp_queue <= #TCQ rdptr_resp_queue + 1;
      if (rd_queue_select_q == REQUEST2_CH)
        rdptr_req2_queue <= #TCQ rdptr_req2_queue + 1;
    end
  end
  generate if (REQ_REORDER) begin: four_queue_rdptr_gen 
    always @(posedge phy_clk) begin
      if (buf_phy_rst_q) begin
        rdptr_req1_queue <= #TCQ 0;
        rdptr_req0_queue <= #TCQ 0;
      end else if (load_backup) begin // backup indication - load backup values
          rdptr_req1_queue <= #TCQ rdptr_backup_req1_queue;
          rdptr_req0_queue <= #TCQ rdptr_backup_req0_queue;
      end else if (rd_tag_ack) begin
        if (rd_queue_select_q == REQUEST1_CH)
          rdptr_req1_queue <= #TCQ rdptr_req1_queue + 1;
        if (rd_queue_select_q == REQUEST0_CH)
          rdptr_req0_queue <= #TCQ rdptr_req0_queue + 1;
      end
    end
  end
  endgenerate

  // update the backup counters whenever we have confirmation that the packet
  // was successfully delivered. After delivery, there is no need to keep
  // that packet any longer. This event occurs subsequent with the clearing
  // of the bit from the Master List.
  reg [4:0] pr_phy_last_ack_q;
  reg [4:0] local_last_acked_q;
  always @(posedge phy_clk) begin
    pr_phy_last_ack_q <= #TCQ PR_phy_last_ack[4:0];
    local_last_acked_q <= #TCQ local_last_acked;
  end

  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      rdptr_backup_resp_queue <= #TCQ 0;
      rdptr_backup_req2_queue <= #TCQ 0;
    end else if (local_last_acked_q != pr_phy_last_ack_q) begin
      if(backup_queue_update == RESPONSE_CH)
        rdptr_backup_resp_queue <= #TCQ rdptr_backup_resp_queue + 1;
      if(backup_queue_update == REQUEST2_CH)
        rdptr_backup_req2_queue <= #TCQ rdptr_backup_req2_queue + 1;
    end
  end

  generate if (REQ_REORDER) begin: four_queue_backup_gen 
    always @(posedge phy_clk) begin
      if (buf_phy_rst_q) begin
        rdptr_backup_req1_queue <= #TCQ 0;
        rdptr_backup_req0_queue <= #TCQ 0;
      end else if (local_last_acked_q != pr_phy_last_ack_q) begin
        if(backup_queue_update == REQUEST1_CH)
          rdptr_backup_req1_queue <= #TCQ rdptr_backup_req1_queue + 1;
        if(backup_queue_update == REQUEST0_CH)
          rdptr_backup_req0_queue <= #TCQ rdptr_backup_req0_queue + 1;
      end
    end
  end
  endgenerate


    // *- ASSERTION (BT_load_backup_and_rd_tag_ack)
    // It is not possible for a backup to occur on the same
    // cycle that an increment indication occurs from the Next Packet Finder.

    // *- COVERAGE (BT_rdptr_resp_queue_enumerate)
    // Enumerate rdptr_resp_queue

    // *- COVERAGE (BT_rdptr_req0_queue_enumerate)
    // Enumerate rdptr_req0_queue

    // *- COVERAGE (BT_rdptr_req1_queue_enumerate)
    // Enumerate rdptr_req1_queue

    // *- COVERAGE (BT_rdptr_req2_queue_enumerate)
    // Enumerate rdptr_req2_queue

    // *- COVERAGE (BT_rdptr_backup_resp_queue_enumerate)
    // Enumerate rdptr_backup_resp_queue

    // *- COVERAGE (BT_rdptr_backup_req0_queue_enumerate)
    // Enumerate rdptr_backup_req0_queue

    // *- COVERAGE (BT_rdptr_backup_req1_queue_enumerate)
    // Enumerate rdptr_backup_req1_queue

    // *- COVERAGE (BT_rdptr_backup_req2_queue_enumerate)
    // Enumerate rdptr_backup_req2_queue

    // *- COVERAGE (BT_rdptr_resp_queue_rollover)
    // Observe rollover on rdptr_resp_queue

    // *- COVERAGE (BT_rdptr_req0_queue_rollover)
    // Observe rollover on rdptr_req0_queue

    // *- COVERAGE (BT_rdptr_req1_queue_rollover)
    // Observe rollover on rdptr_req1_queue

    // *- COVERAGE (BT_rdptr_req2_queue_rollover)
    // Observe rollover on rdptr_req2_queue

    // *- COVERAGE (BT_rdptr_backup_resp_queue_rollover)
    // Observe rollover on rdptr_backup_resp_queue

    // *- COVERAGE (BT_rdptr_backup_req0_queue_rollover)
    // Observe rollover on rdptr_backup_req0_queue

    // *- COVERAGE (BT_rdptr_backup_req1_queue_rollover)
    // Observe rollover on rdptr_backup_req1_queue

    // *- COVERAGE (BT_rdptr_backup_req2_queue_rollover)
    // Observe rollover on rdptr_backup_req2_queue

    // *- ASSERTION (BT_rdptr_queue_increment)
    // It is only possible for one rdptr_*_queue counter to increment at a time.

    // *- ASSERTION (BT_rdptr_backup_queue_increment)
    // It is only possible for one rdptr_backup_*_queue counter to increment at a time.

    // *- COVERAGE (BT_rdptr_queue_cross_rdptr_backup_queue)
    // Cross load_backup with each rdptr_*_queue, crossed with
    // rdptr_backup_*_queue, crossed with TX_DEPTH
    // Interesting values of the queue counters: 0, 1, 2, ...,
    // TX_DEPTH-2, TX_DEPTH-1, TX_DEPTH

    // *- ASSERTION (BT_resp_backup_passes_rdptr)
    // It is not possible for backup_resp_queue counter to pass resp_queue

    // *- ASSERTION (BT_req0_backup_passes_rdptr)
    // It is not possible for backup_req0_queue counter to pass req0_queue

    // *- ASSERTION (BT_req1_backup_passes_rdptr)
    // It is not possible for backup_req1_queue counter to pass req1_queue

    // *- ASSERTION (BT_req2_backup_passes_rdptr)
    // It is not possible for backup_req2_queue counter to pass req2_queue

  // }}} end Read Pointer Maintenance --


  // {{{ Next Packet Finder ---------

  // Need a simple way to determine if there is a packet pending in one of the
  // queues. If the values of the counters are not equal, then there is a packet pending.
  wire       resp_pending = !(wrptr_resp_queue == rdptr_resp_queue);
  wire       req2_pending = !(wrptr_req2_queue == rdptr_req2_queue);
    // These two removed when REQ_REORDER = 0
  wire       req1_pending = !(wrptr_req1_queue == rdptr_req1_queue);
  wire       req0_pending = !(wrptr_req0_queue == rdptr_req0_queue);

  wire       resp_prio_mask;
  wire       prio2_mask, prio1_mask, prio0_mask;
  reg        prio2_mask_q, prio1_mask_q, prio0_mask_q;


  // Generate the signal that determines flow control. This will be sent on to the PHY OLLM RX.
  generate if (RX_FC_ONLY || !REQ_REORDER) begin: rx_fc_only_gen
    always @* begin
      // in order to synthesize in xst, there must be at least one item in the sensitivity list.
      if (buf_phy_rst_q)
        BT_tx_flow_control = 1'b0;
      else
        BT_tx_flow_control = 1'b0;
    end
  end else                 begin: rxtx_fc_gen
    always @(posedge phy_clk) begin
      if (buf_phy_rst_q)
        BT_tx_flow_control <= #TCQ 1'b1;
      else if (BC_force_rx_flow)
        BT_tx_flow_control <= #TCQ 1'b0;
      else
        BT_tx_flow_control <= #TCQ ~&PR_phy_rcvd_buf_stat;
    end
  end
  endgenerate


  // When in Transmitter Flow control (tbuf_stat != 'hFF), mask pending
  // packets based on the values of the watermarks. Otherwise, there are no masks.
  generate if (!RX_FC_ONLY) begin: rxtx_mask_gen
    assign     resp_prio_mask = (link_free_buffer != 0)             || !BT_tx_flow_control;
    assign     prio2_mask     = (link_free_buffer >= BC_watermark2) || !BT_tx_flow_control;
    assign     prio1_mask     = (link_free_buffer >= BC_watermark1) || !BT_tx_flow_control;
    assign     prio0_mask     = (link_free_buffer >= BC_watermark0) || !BT_tx_flow_control;
  end else                  begin: rx_only_mask_gen
    assign     resp_prio_mask = 1'b1;
    assign     prio2_mask     = 1'b1;
    assign     prio1_mask     = 1'b1;
    assign     prio0_mask     = 1'b1;
  end
  endgenerate
  generate if (!RX_FC_ONLY) begin: prio_mask_q_gen
    always @(posedge phy_clk) begin
      if (rd_tag_ack_d) begin
        prio2_mask_q <= #TCQ prio2_mask;
        prio1_mask_q <= #TCQ prio1_mask;
        prio0_mask_q <= #TCQ prio0_mask;
      end
    end
  end else                  begin: fake_prio_mask_q_gen
    always @(posedge phy_clk) begin
      prio2_mask_q <= #TCQ 1'b1;
      prio1_mask_q <= #TCQ 1'b1;
      prio0_mask_q <= #TCQ 1'b1;
    end
  end
  endgenerate


  // final accumulation for the list of pending packets by queue.
  generate if (REQ_REORDER) begin: four_queue_pending_list_gen 
    assign raw_pending_list = {resp_pending, req2_pending, req1_pending, req0_pending};
    assign pending_list     = {resp_pending && resp_prio_mask,
                               req2_pending && prio2_mask,
                               req1_pending && prio1_mask,
                               req0_pending && prio0_mask};
  end else                  begin: two_queue_pending_list_gen
    assign raw_pending_list = {resp_pending, req2_pending, 1'b0, 1'b0};
    assign pending_list     = {resp_pending && resp_prio_mask,
                               req2_pending && prio2_mask,
                               1'b0,
                               1'b0};
  end
  endgenerate


  // this is a priority based evaluation. Regardless of the status of a lower
  // priority, a higher priority gets selected.
  always @* begin
    casex (raw_pending_list)
      // in order of priority, highest to lowest
      4'b1xxx : rd_queue_select = RESPONSE_CH;
      4'b01xx : rd_queue_select = REQUEST2_CH;
      4'b001x : rd_queue_select = REQUEST1_CH;
      4'b0001 : rd_queue_select = REQUEST0_CH;
      default : rd_queue_select = 'hx;
    endcase
  end
  // register the select to the mux. We'll use this to remember which address
  // we sent to the Read Port Controller. This is important when the select
  // line changes near the time when the read controller starts a new packet.
  always @(posedge phy_clk) begin
    if (rd_tag_ack_d)
      rd_queue_select_q <= #TCQ rd_queue_select;
  end


  // qualify the address tag to the Read Port Controller by indicating if it
  // is valid. If it being acked on the current cycle, release valid,
  // otherwise, it will appear to be a new address to the read address logic.
  // NOTE - we compare next_fm and last_ack to make sure we don't transmit more than 31 packets.
  // There is nothing that prevents us from transmitting all 32 packets, except that there
  // is no way to differentiate between a PNA with no implicit ACKs and a PNA with an inplicit ACK of 32
  // packets. In both cases, the last_ack value will match. So, we avoid the whole situation by only
  // allowing 31 outstanding packets (found by comparing these two values).
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      rd_tag_valid <= #TCQ 1'b0;
    else
      rd_tag_valid <= #TCQ (|pending_list) && (PR_phy_rcvd_buf_stat != free_buf_partial_sum) &&
                            &transmit_enable && !load_backup_d &&
                            // following lines prevent more than 31 packets being outstanding
                            (PR_phy_last_ack[4:0] != local_next_acked[4:0]);
// FIXME - CFR - remove once regressions pass successfully
//                            (PR_phy_last_ack[4:0] != PT_phy_next_fm[4:0]) &&
//                            (PR_phy_last_ack[4:0] != (PT_phy_next_fm[4:0] + 5'h1));
  end


  // corner-case protection logic- Specifically for TX flow control, because
  // of the latency between some paths, an occasional request may pass through
  // just as a response is getting ready. If the watermarks are changing at
  // the same time, we may accidentally bump the request's priority because we
  // think it is a response. This logic prevents this very rare occurrance.
  always @(posedge phy_clk) begin
    if (rd_tag_ack_pulse)
      transmitting_resp <= #TCQ rd_queue_select_q == RESPONSE_CH;
  end


  // When in Transmitter Controlled Flow Control, the logic must evaluate how
  // many free locations exist in the link partner's buffer. The link partner
  // provides this information with PR_phy_rcvd_buf_stat. However, there are also
  // packets that have not been accounted for. Those packets may be
  // quantified by subtracting the difference between PR_phy_last_ack and
  // PT_phy_next_fm.
  // For the partial sum, note when there are no outstanding packets, the
  // difference is actually 1. i.e. next = 1, last = 0; this means there are
  // no outstanding packets. So, subtract 1 from next.
  assign free_buf_partial_sum = local_next_acked - PR_phy_last_ack[4:0] - 1;

  // The number of free buffer locations in the link partner becomes the
  // difference.
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      link_free_buffer <= #TCQ 6'h3F;
    else if (((PR_phy_rcvd_buf_stat > ({1'b0, free_buf_partial_sum} + C_TX_FC_TUNER)) ||
              (free_buf_partial_sum == 0)) &&
             (local_next_acked != PR_phy_last_ack[4:0]))
      link_free_buffer <= #TCQ PR_phy_rcvd_buf_stat - {1'b0, free_buf_partial_sum} - C_TX_FC_TUNER;
    else
      link_free_buffer <= #TCQ 6'h0;
  end


  // TX flow control priority adjust -
  // This logic is used in the case of TX flow control. It jumps directly to
  // the proper priority for responses.
  // Only generate if we are not in forced Receiver flow control.
  generate if (!RX_FC_ONLY) begin: tx_prio_gen
    always @* begin
      casex ({prio2_mask_q, prio1_mask_q, prio0_mask_q})
        3'b111  : tx_prio_adjust =  2'h0;
        3'b110  : tx_prio_adjust =  2'h1;
        3'b100  : tx_prio_adjust =  2'h2;
        3'b000  : tx_prio_adjust =  2'h3;
        default : tx_prio_adjust =  2'hx;
      endcase
    end
  end
  endgenerate


    // *- ASSERTION (BT_bram_raddr_u_is_x)
    // There will never be a time when bram_raddr_u is X when there is a read.

    // *- ASSERTION (BT_link_free_buffer_underrun)
    // link_free_buffer can only arrive at 0 from either 0 or 1. i.e.
    // We should never see link_free_buffer underrun: (high-value -> 00)

    // *- COVERAGE (BT_link_free_buffer_enumerate)
    // Enumerate link_free_buffer

    // *- COVERAGE (BT_pending_list_enumerate)
    // Enumerate pending_list

    // *- COVERAGE (BT_link_free_buffer_cross_pending)
    // Cross all *_pending signals with link_free_buffer = {0, 1, 2, 3, 4+}

    // *- COVERAGE (BT_pending_cross_masks)
    // Cross all *_pending signals with the masks

    // *- COVERAGE (BT_free_buf_partial_sum_cross_rewind)
    // Cross free_buf_partial_sum with PT_phy_rewind

  // }}} end Next Packet Finder -----


  // {{{ Address Select -------------

  // mux the tags coming from the distributed memory, resulting in the next
  // read tag location.
  generate if (REQ_REORDER) begin: four_queue_next_read_tag_gen
    always @* begin
      case (rd_queue_select)
        // in order of priority, highest to lowest
        RESPONSE_CH : next_read_tag = rs_read_tag;
        REQUEST2_CH : next_read_tag = r2_read_tag;
        REQUEST1_CH : next_read_tag = r1_read_tag;
        REQUEST0_CH : next_read_tag = r0_read_tag;
        default     : next_read_tag = 'hx;
      endcase
    end
  end else                  begin: two_queue_next_read_tag_gen
    always @* begin
      case (rd_queue_select)
        // in order of priority, highest to lowest
        RESPONSE_CH : next_read_tag = rs_read_tag;
        REQUEST2_CH : next_read_tag = r2_read_tag;
        default     : next_read_tag = 'hx;
      endcase
    end
  end
  endgenerate
  // }}} end Address Select ---------


  // {{{ Read Port Controller -------
  reg    bt_bram_rd_frame, bt_bram_rd_frame_q; // asserted while in a packet
  reg    update_window, update_window_q;       // asserted while outside of a packet
  reg    set_update_window;

  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      bt_bram_rd_frame_q <= #TCQ 1'b0;
      update_window_q    <= #TCQ 1'b1;
      rd_tag_ack_pulse   <= #TCQ 1'b0;
    end else begin
      bt_bram_rd_frame_q <= #TCQ bt_bram_rd_frame;
      update_window_q    <= #TCQ update_window;
      rd_tag_ack_pulse   <= #TCQ rd_tag_ack_d;
    end
  end

  // generate a signal to acknowledge which tag queue we'll be pulling from and to stop all
  // deliberation towards reordering.
  always @* begin
    update_window = update_window_q;
    // clear two cycles before TSTART for multi-cycle packets
    if (rd_tag_ack_pulse && !PT_phy_rewind)
      update_window = 1'b0;
    else if (set_update_window)
      update_window = 1'b1;
  end
  always @* begin
    set_update_window = 1'b0;
    // always allow an update on single cycle packets
    // for multi-cycle packets, wait for the next-to-last phase
    if (btb_tx_last && PT_phyt_tready && (BT_phyt_tvalid || bt_phyt_tvalid_d[1]))
      set_update_window = 1'b1;
    // for small packets that are fewer cycles than the depth of the pipeline
    else if (btb_tx_last && !BT_phyt_tvalid)
      set_update_window = 1'b1;
    // finally, this is a reset upon rewind
    else if (PT_phy_rewind)
      set_update_window = 1'b1;
  end


  // create the acknowledgement signal when the logic captures the next_read_tag.
  assign rd_tag_ack_d = |pending_list && rd_tag_valid && update_window && &transmit_enable && bt_phyt_advance;
  assign rd_tag_ack   = rd_tag_ack_hold && bt_phyt_advance;

  // simply registering rd_tag_ack_d is not sufficient to determine if we can
  // move to the next packet. This is true in the case where TREADY deasserts
  // on the very last data phase of the previous packet (when TLAST is asserted).
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      rd_tag_ack_hold <= #TCQ 1'b0;
    end else begin
      rd_tag_ack_hold <= #TCQ rd_tag_ack_d || (rd_tag_ack_hold && !bt_phyt_advance && !PT_phy_rewind);
    end
  end


  // Read enable generation -
  // only read during an active packet. This specifically prevents old eof
  // signals from interfereing with the new packet.
  // Create a frame signal which indicates when it's safe to read from the memory.
  // It is safe to read from memory so long as tags keep getting acknowledged
  always @* begin
    bt_bram_rd_frame = bt_bram_rd_frame_q;
    // set upon acking the tag
    if (rd_tag_ack && !PT_phy_rewind)
      bt_bram_rd_frame = 1'b1;
    else if (set_update_window)
      bt_bram_rd_frame = 1'b0;
  end
  assign bt_bram_rd = bt_bram_rd_frame && bt_phyt_advance;


  // Read address generation -
  // The lower portion of the address resets to zero. It also loads zero when
  // EOF is observed. Otherwise, it incrments by one every time valid data is present.
  // The upper portion of the address loads from the Address Select only when
  // it has completed the previous transaction.
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      bram_raddr_u <= #TCQ 0;
    end else if (rd_tag_valid && update_window) begin
      bram_raddr_u <= #TCQ next_read_tag;
    end
  end
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      bram_raddr_l <= #TCQ 0;
    end else if (bt_bram_rd) begin
      bram_raddr_l <= #TCQ bram_raddr_l + 1;
    end else if (set_update_window) begin
      bram_raddr_l <= #TCQ 0;
    end
  end


    // *- COVERAGE (BT_bt_bram_rd_two_after_tlast)
    // Observe a read two cycles after tlast asserts from an address whose lower bits are zero
    // Between cycles, observe that bt_bram_rd is low - i.e. observe a gap of 2 cycles between packets

    // *- COVERAGE (BT_bt_bram_rd_three_after_tlast)
    // Observe a read three cycles after tlast asserts from an address whose lower bits are zero
    // Between cycles, observe that bt_bram_rd is low - i.e. observe a gap of 3 cycles between packets

    // *- COVERAGE (BT_bt_bram_rd_four_after_tlast)
    // Observe a read four cycles after tlast asserts from an address whose lower bits are zero
    // Between cycles, observe that bt_bram_rd is low

    // *- COVERAGE (BT_bt_bram_raddr_non_zero_reset)
    // Observe a reset when both the upper and lower portions of the read address are non-zero

    // *- COVERAGE (BT_bram_raddr_non_zero_reset)
    // Observe a reset when both the upper and lower portions of the read address are non-zero

    // *- ASSERTION (BT_rd_tag_ack_d_and_rewind)
    // It is not possible for rd_tag_ack_d to assert on the same cycle as a rewind

    // *- ASSERTION (BT_rd_tag_ack_d_and_rewind_minus_one)
    // It is not possible for rd_tag_ack_d to assert one cycle after a rewind

    // *- ASSERTION (BT_rd_tag_ack_d_and_rewind_minus_two)
    // It is not possible for rd_tag_ack_d to assert two cycles after a rewind

    // *- COVERAGE (BT_rd_tag_ack_d_and_rewind_plus_one)
    // Observe rewind asserted one cycle after rd_tag_ack_d

    // *- COVERAGE (BT_rd_tag_ack_d_and_rewind_plus_two)
    // Observe rewind asserted two cycles after rd_tag_ack_d

  // }}} end Read Port Controller ---


  // {{{ ACK ID Maintenance ---------

  reg                  load_backup_q;
  reg  [4:0]           local_next_acked_q, local_next_acked_qq;
  reg  [C_TAG_LEN-1:0] next_read_tag_q, next_read_tag_qq;
  reg  [1:0]           rd_queue_select_qq;
  reg  [1:0]           observed_rewind_already;

  // declare the memories implicitly. There are 32 possible storage locations,
  // so we must keep locations for all of them. One of these memories holds
  // tag information while the other holds queue information. Popping each one
  // off causes the removal of that tag from record.
  //
  // initialize queue_lookup to be something other than the response channel
  // lest we accidentally bump priority when we shouldn't.
  (* ram_style = "distributed" *)
  reg  [C_TAG_LEN-1:0] tag_lookup   [0:31];
  (* ram_style = "distributed" *)
  reg  [1:0]           queue_lookup [0:31];
  integer ii, jj;

// added below macro to fix the CR# 735137
// synthesis translate_off 
  initial for (ii = 0; ii < 32; ii = ii + 1) tag_lookup[ii] = 0;
  initial for (jj = 0; jj < 32; jj = jj + 1) queue_lookup[jj] = REQUEST0_CH;
// synthesis translate_on


  // generate the read address into the dist ram. This is used to index
  // into both the queue lookup and the tag lookup.
  // Why is load_backup used here? Whenever there is a rewind, we have to
  // grab the queue and tag information of the retried packet in order to
  // know if we need to bump priority or not.
  wire [4:0] ack_tag_rd_addr = load_backup ? PT_phy_next_fm[4:0] : local_last_acked;


  // local copies of PR_phy_last_ack and PT_phy_next_fm - renamed to more
  // comprehendable names.
  // generate local next ack id logic. The value in this counter should lead
  // the real next ack id (tnext_fm) by a few cycles. We'll use this to write
  // information into the distributed ram. The ack id always increments by
  // one unless there is a retry condition. In that case, the link partner
  // tells us where to start up again.
  // The delay version is used specifically for determining if there are no
  // outstanding packets to bump a priority on. We cannot use the regular
  // count version because it increments before we are certain that the packet
  // has been sent.
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      local_next_acked       <= #TCQ 5'h0;
      local_next_acked_delay <= #TCQ 5'h0;
    // don't increment if we see a rewind 
    end else begin
      if (BT_phyt_tlast && BT_phyt_tvalid && PT_phyt_tready) begin
        local_next_acked_delay <= #TCQ local_next_acked_delay + 1;
      // unfortunately, we have to do this in order to get the local value to be
      // accurate against the external value. This is important because the PHY
      // can NAK a packet that has already been ACKed. This is a special case
      // that we must consider.
      end else if (load_backup) begin
        local_next_acked_delay <= #TCQ PT_phy_next_fm[4:0];
      end

      if (rd_tag_ack && !PT_phy_rewind) begin
        local_next_acked <= #TCQ local_next_acked + 1;
      // unfortunately, we have to do this in order to get the local value to be
      // accurate against the external value. This is important because the PHY
      // can NAK a packet that has already been ACKed. This is a special case
      // that we must consider.
      end else if (load_backup) begin
        local_next_acked <= #TCQ PT_phy_next_fm[4:0];
      end
    end
  end



  // unfortunate requirement - we can witness back-to-back rewinds. So,
  // while we're handling the first one, a second one can come and hose up how
  // we're handling the first discontinue. So, we must wait to actually place
  // the pointers and tag information into the dist ram until we witness
  // a real assertion of sof.
  // when we witness rd_tag_ack_d, store pointers into memory, as well as the
  // values. If we could ensure that back-to-back discontinues would not
  // occur, we would store directly into memory upon the assertion of
  // rd_tag_ack_d.
  always @(posedge phy_clk) begin
    if (rd_tag_ack_d) begin
      local_next_acked_q <= #TCQ local_next_acked;
      next_read_tag_q    <= #TCQ next_read_tag;
    end
  end
  always @(posedge phy_clk) begin
    local_next_acked_qq <= #TCQ local_next_acked_q;
    next_read_tag_qq    <= #TCQ next_read_tag_q;
    rd_queue_select_qq  <= #TCQ rd_queue_select_q;
  end


  // generate the local last ack id logic. Everytime the PHY layer updates
  // the last ack signal, we follow suit. The result is that we pop off a tag
  // reference from the tag lookup and a queue reference from the queue lookup.
  assign bt_packet_ack = (local_last_acked != PR_phy_last_ack[4:0]);
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      bt_packet_ack_q  <= #TCQ 1'b0;
      local_last_acked <= #TCQ 5'h1F;
    end else begin
      bt_packet_ack_q  <= #TCQ bt_packet_ack;
      if (bt_packet_ack) begin
        local_last_acked <= #TCQ local_last_acked + 1;
      end
    end
  end


  // read-side operation-
  // keep this clean to ensure the we get the structure we actually want.
  // The output of this memory is used to clear the master list when a packet
  // finally gets acknowledged. Also, it is used when bumping a priority.
  assign current_ack_tag_d = tag_lookup[ack_tag_rd_addr];


  // write-side operation-
  // Store the next read tag for the sole purpose of if it gets retried at a later date.
  // Why are we using _qq for address and write value?
  // The first stage (_q) values are captured on the very cycle that we determine which queue to pick from.
  // The second stage (_qq) is required because a second transfer can start before we record the first transfer.
  // keep this clean to ensure the we get the structure we actually want.
  always @(posedge phy_clk) begin
    if (bt_phyt_tstart)
      tag_lookup[local_next_acked_qq] <= #TCQ next_read_tag_qq;
  end


  // generate the distributed tag for the acknowledged packet.
  always @(posedge phy_clk) begin
    current_ack_tag <= #TCQ current_ack_tag_d;
  end


  // backup counter increment -
  // generate the queue reference signals associated with the backup counters.
  // Whenever a packet gets acked, send the appropriate increment signal.
  // This is the sole purpose of the queue lookup memory.
  // Why are we using _qq for address and write value?
  // The first stage (_q) values are captured on the very cycle that we determine which queue to pick from.
  // The second stage (_qq) is required because a second transfer can start before we record the first transfer.
  // keep this clean to ensure the we get the structure we actually want.
  always @(posedge phy_clk) begin
    if (bt_phyt_tstart)
      queue_lookup[local_next_acked_qq] <= #TCQ rd_queue_select_qq;
  end


  // keep this clean to ensure the we get the structure we actually want.
  // read operation
  assign backup_queue_update = queue_lookup[ack_tag_rd_addr];


  // generate transmit enable-
  // The only time this module interferes with operation is when things must
  // back up. In that case, the transmit enable signal prevents any further
  // packets from being transmitted until the pointers have all been backed up.
  reg  eval_for_backup, eval_for_backup_q;
  wire set_load_backup_d;
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      load_backup        <= #TCQ 1'b0;
      load_backup_q      <= #TCQ 1'b0;
      transmit_enable[1] <= #TCQ 1'b1;
      pr_phy_rewind_q    <= #TCQ 1'b0;
      eval_for_backup_q  <= #TCQ 1'b0;
    end else begin
      load_backup        <= #TCQ load_backup_d;
      load_backup_q      <= #TCQ load_backup;
      transmit_enable[1] <= #TCQ transmit_enable[0];
      pr_phy_rewind_q    <= #TCQ PT_phy_rewind;
      eval_for_backup_q  <= #TCQ eval_for_backup;
    end
  end
  always @* begin
    if (PT_phy_rewind)
      transmit_enable[0] = 1'b0;
    else if (load_backup_q && !PT_phy_rewind && !pr_phy_rewind_q)
      transmit_enable[0] = 1'b1;
    else
      transmit_enable[0] = transmit_enable[1];
  end


  // kickoff the recovery process. Once all acked packets have been cleared,
  // it should take only 4 cycles to start resending packets again.
  always @* begin
    eval_for_backup = eval_for_backup_q;
    if (!PT_phy_rewind && pr_phy_rewind_q)
      eval_for_backup = 1'b1;
    else if (load_backup_d)
      eval_for_backup = 1'b0;
  end
  assign set_load_backup_d = eval_for_backup && (local_last_acked == PR_phy_last_ack[4:0]) &&
                             !(load_backup_d || load_backup);
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      load_backup_d <= #TCQ 1'b0;
    else if (set_load_backup_d)
      load_backup_d <= #TCQ 1'b1;
    else
      load_backup_d <= #TCQ 1'b0;
  end

  // qualifies whether the Priority Adjust actually needs to take action.
  // a rewind can happen on an empty buffer. You can usually see that
  // when next_acked and next_fm are not equal. However, a completey full
  // and completely empty buffer look the same. For that reason, we do not allow all 32
  // packets to be outstanding.
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      resp_retry <= #TCQ 1'b0;
    else if (load_backup && (local_next_acked_delay != PT_phy_next_fm[4:0]))
      resp_retry <= #TCQ backup_queue_update == RESPONSE_CH;
    else if (load_backup && (local_next_acked_delay == PT_phy_next_fm[4:0]) && !observed_rewind_already[1])
      resp_retry <= #TCQ 1'b0;
    else if (!alt_prio_available && alt_prio_available_q)
      resp_retry <= #TCQ 1'b0;
  end
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      observed_rewind_already <= #TCQ 2'b0;
    else if (!PT_phy_rewind && pr_phy_rewind_q)
      observed_rewind_already <= #TCQ {observed_rewind_already[0], 1'b1};
    else if (bt_phyt_tstart && PT_phyt_tready && !PT_phy_rewind)
      observed_rewind_already <= #TCQ 2'b0;
  end


    // *- COVERAGE (BT_local_next_acked_enumerate)
    // Enumerate local_next_acked

    // *- COVERAGE (BT_local_next_acked_rollover)
    // Observe local_next_acked rolls over

    // *- COVERAGE (BT_local_last_acked_enumerate)
    // Enumerate local_last_acked

    // *- COVERAGE (BT_local_last_acked_rollover)
    // Observe local_last_acked rolls over

    // *- COVERAGE (BT_local_next_acked_cross_pt_phy_next_fm)
    // Cover next_fm = PT_phy_next_fm, PT_phy_next_fm+1, PT_phy_next_fm+2

    // *- ASSERTION (BT_local_next_acked_behavior)
    // Except on rewind, local_next_acked may not be any value other than
    // PT_phy_next_fm, PT_phy_next_fm+1, or PT_phy_next_fm+2

    // *- COVERAGE (BT_bt_phyt_tstart_and_rewind)
    // Observe rewind asserted on the same cycle as bt_phyt_tstart

    // *- ASSERTION (BT_bt_phyt_tstart_and_rewind_minus_one)
    // It is not possible for bt_phyt_tstart to assert one cycle after a rewind

    // *- ASSERTION (BT_bt_phyt_tstart_and_rewind_minus_two)
    // It is not possible for bt_phyt_tstart to assert two cycles after a rewind

    // *- COVERAGE (BT_bt_phyt_tstart_and_rewind_plus_one)
    // Observe rewind asserted one cycle after bt_phyt_tstart

    // *- COVERAGE (BT_bt_phyt_tstart_and_rewind_plus_two)
    // Observe rewind asserted two cycles after bt_phyt_tstart

  // }}} end ACK ID Maintenance -----


  // {{{ Control Signal Drivers -----

  // generate the advance signal -
  // Indicates when to push data from the bram or pull from the interface through the pipeline
  assign bt_phyt_advance = PT_phyt_tready || !BT_phyt_tvalid;


  // generate TSTART -
  // This is signal is mocked to look like the AXI interface. While it is
  // not used in the interface, it is a very useful signal internally.
  // Indicates the first data beat of a packet.
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      bt_phyt_tstart <= #TCQ 1'b0;
    else if (PT_phy_rewind)
      bt_phyt_tstart <= #TCQ 1'b0;
    else if (bt_phyt_advance)
      bt_phyt_tstart <= #TCQ btb_tx_start;
  end


  // generate TLAST -
  // generally forward the TLAST from the block ram. However, upon
  // a discontinue, issue a TLAST on the next cycle, assuming there was not a
  // TLAST on the previous cycle.
  reg  bt_phyt_src_dsc, bt_phyt_src_dsc_q;
  always @* begin
    if (PT_phy_rewind && bt_phyt_tvalid_d[1]) // Set src_dsc when in mid packet
      bt_phyt_src_dsc = 1'b1;
    else if (BT_phyt_tuser[0]) // Clear src_dsc any time the interface advances
      bt_phyt_src_dsc = 1'b0;
    else
      bt_phyt_src_dsc = bt_phyt_src_dsc_q;
  end
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      bt_phyt_src_dsc_q <= #TCQ 1'b0;
    else
      bt_phyt_src_dsc_q <= #TCQ bt_phyt_src_dsc;
  end

  assign bt_phyt_tlast_d = btb_tx_last || bt_phyt_src_dsc;
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      BT_phyt_tlast <= #TCQ 1'b0;
    end else if (bt_phyt_advance) begin
      BT_phyt_tlast <= #TCQ bt_phyt_tlast_d && bt_phyt_tvalid_d[1];
    end
  end


  // generate TUSER -
  // Just pass along from the BRAM
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      BT_phyt_tuser <= #TCQ 8'h0;
    else if (bt_phyt_advance)
      BT_phyt_tuser <= #TCQ {5'h0, btb_tx_user, bt_phyt_src_dsc};
  end



  // generate TVALID -
  // never assert ready outside of a packet. always have it asserted during
  // a packet. This signal carries forward and is pipelined to match the 
  // path that the data travels. Since there are three stages of pipeline,
  // there are three stages of the valid signal. It is important that this
  // travel along with the data in order to know how to handle the data.
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      bt_phyt_tvalid_d[0] <= #TCQ 1'b0;
    end else if (PT_phy_rewind) begin
      bt_phyt_tvalid_d[0] <= #TCQ 1'b0;
    end else if (bt_bram_rd) begin
      if (btb_tx_bram_last && (bt_bram_raddr[C_INDEX_LEN-1:0] != 0)) begin
        bt_phyt_tvalid_d[0] <= #TCQ 1'b0;
      end else begin
        bt_phyt_tvalid_d[0] <= #TCQ 1'b1;
      end
    end else if (bt_phyt_advance) begin
      bt_phyt_tvalid_d[0] <= #TCQ 1'b0;
    end
  end
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      bt_phyt_tvalid_d[1] <= #TCQ 1'b0;
      BT_phyt_tvalid      <= #TCQ 1'b0;
    end else if (bt_phyt_advance) begin
      bt_phyt_tvalid_d[1] <= #TCQ bt_phyt_tvalid_d[0] && !PT_phy_rewind;
      BT_phyt_tvalid      <= #TCQ bt_phyt_tvalid_d[1] && !(PT_phy_rewind && !BT_phyt_tvalid);
    end
  end


  // generate TSTRB -
  // Reconstruct the strobe. 
  // When not in a packet, strobe = 00
  // When in a packet and not the last cycle, strobe = FF
  // When on the last cycle, expand the strobe from the BRAM
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      BT_phyt_tkeep <= #TCQ 8'h0;
    end else if (bt_phyt_advance) begin
      if (!bt_phyt_tvalid_d[1]) begin
        BT_phyt_tkeep <= #TCQ 8'h0;
      end else if (!bt_phyt_tlast_d) begin
        BT_phyt_tkeep <= #TCQ 8'hFF;
      end else begin
        BT_phyt_tkeep <= #TCQ {1'b0, btb_tx_keep[2], btb_tx_keep[2], btb_tx_keep[1], 
                               btb_tx_keep[1], btb_tx_keep[0], btb_tx_keep[0], 1'b1};
      end
    end
  end


  // generate TDATA -
  // For the most part, data comes directly from Block RAM. This logic MUXs
  // in alternate priorities when required.
  wire [1:0]           existing_priority = btb_tx_data[7:6];
  reg  [C_TAG_LEN-1:0] bram_raddr_u_q;
  wire                 adjust_with_rx_prio = // mux condition to take adjusted rx priority
                        btb_tx_start && alt_prio_available && (bram_raddr_u_q == tag_marker);
  wire                 adjust_with_tx_prio = // mux condition to take adjusted tx priority
                        btb_tx_start && transmitting_resp && (tx_prio_adjust > existing_priority);
  wire                 tx_is_greater_than_rx_prio = // used to determine which prio to take
                        transmitting_resp && (tx_prio_adjust > existing_priority && tx_prio_adjust > rx_prio_adjust);

  generate if (!RX_FC_ONLY) begin: rxtx_priority_gen
    always @(posedge phy_clk) begin
      // RX flow control option for bumping priority
      // increment by one until acceptance.
      if (buf_phy_rst_q) begin
        BT_phyt_tdata <= #TCQ 64'h0;
      end else if (bt_phyt_advance) begin
        // is the tx bump higher and valid? If so, skip to next condition
        if (adjust_with_rx_prio && !tx_is_greater_than_rx_prio) begin
          BT_phyt_tdata <= #TCQ {btb_tx_data[63:8], rx_prio_adjust, btb_tx_data[5:0]};
        // TX flow control option for bumping priority - immediate increment to the proper value.
        end else if (adjust_with_tx_prio) begin
          BT_phyt_tdata <= #TCQ {btb_tx_data[63:8], tx_prio_adjust, btb_tx_data[5:0]};
        end else begin // standard procedure
          BT_phyt_tdata <= #TCQ btb_tx_data;
        end 
      end
    end

  end else                  begin: rx_only_priority_gen
    always @(posedge phy_clk) begin
      if (buf_phy_rst_q) begin
        BT_phyt_tdata <= #TCQ 64'h0;
      end else if (bt_phyt_advance) begin
        // RX flow control option for bumping priority - increment by one until acceptance.
        if (adjust_with_rx_prio) begin
          BT_phyt_tdata <= #TCQ {btb_tx_data[63:8], rx_prio_adjust, btb_tx_data[5:0]};
        end else begin // standard procedure
          BT_phyt_tdata <= #TCQ btb_tx_data;
        end
      end
    end

  end
  endgenerate

  always @(posedge phy_clk) begin
    if (bt_phyt_advance)
      bram_raddr_u_q <= #TCQ bram_raddr_u;
  end


    // *- COVERAGE (BT_rewind_on_tlast)
    // Observe PHY asserts rewind on the last cycle of a transaction, the
    // same cycle when TLAST is asserted.

    // *- COVERAGE (BT_rewind_one_after_tlast)
    // Observe PHY asserts rewind one cycle after the last cycle of a transaction.

    // *- COVERAGE (BT_rewind_two_after_tlast)
    // Observe PHY asserts rewind two cycles after the last cycle of a transaction.

    // *- COVERAGE (BT_rewind_on_start)
    // Observe PHY asserts rewind on the same cycle as the first data beat of a packet.

    // *- COVERAGE (BT_rewind_on_second_beat)
    // Observe PHY asserts rewind on the second cycle of a packet.

    // *- COVERAGE (BT_rewind_before_start)
    // Observe PHY asserts rewind one cycle before the first data beat of a packet.

    // *- COVERAGE (BT_rewind_single_cycle)
    // Observe a rewind asserted for only one cycle

    // *- COVERAGE (BT_rewind_multi_cycle)
    // Observe a rewind asserted for 8 or more cycles

    // *- COVERAGE (BT_rewind_repeat)
    // Observe consecutive assertions of rewind, without the beginning of a new packet between them.

  // }}} end Control Signal Drivers -

endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/buf/buf_cfg/srio_gen2_v4_1_16_buf_cfg_top.v#1 $
//----------------------------------------------------------------------
//
// BUF_CFG_TOP
// Description:
// This module contains the configuration registers for the Buffer.
//
// It uses an AXI-Lite interface to the Configuration Fabric, and has a
// BUF core interface for transfer of control and status information.
//
// No clock relationship between cfg_clk and phy_clk is assumed.
//
// Hierarchy:
// BUF_TOP
//    |______BUF_CFG_TOP <-- this module
//              |______CFG_AXI (in hdl/common/)
//              |______BUF_CFG_REG
// ---------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)

module srio_gen2_v4_1_16_buf_cfg_top
  #(
    parameter TCQ         = 100,
    parameter TX_DEPTH    = 32,   // TX buffer depth {8, 16, 32}
    parameter RX_DEPTH    = 32,   // RX buffer depth {8, 16, 32}
    parameter RX_FC_ONLY  = 0,    // RX Flow Control Only {0, 1}
    parameter UNIFIED_CLK = 0,    // phy_clk = log_clk {0, 1}
    parameter REQ_REORDER = 1,    // Request reordering enabled {0, 1}
    parameter WM0         = 3,    // Watermark 0 reset value {WM0 < 64}
    parameter WM1         = 2,    // Watermark 1 reset value {WM0 > WM1 > WM2}
    parameter WM2         = 1,    // Watermark 2 reset value {WM2 > 0}
    parameter IDLE2       = 0)    // IDLE2 sequence support
  (
    // {{{ Port Declarations ---------------
    // System Signals
    input             phy_clk,                // PHY interface clock
    input             buf_phy_rst,            // Reset for PHY clock domain
    input             cfg_clk,                // CFG Interface user clock
    input             cfg_rst,                // Reset for CFG clk domain

    // Buffer Interface
    input             BT_tx_flow_control,     // TX Flow Control Mode
    input             PP_idle2_selected,      // OPLM has trained to use IDLE2 sequence
    output     [5:0]  BC_watermark0,          // Watermark 0
    output     [5:0]  BC_watermark1,          // Watermark 1
    output     [5:0]  BC_watermark2,          // Watermark 2
    output            BC_force_rx_flow,       // Force the Buffer into RX Flow Control mode

    // Configuration Fabric Interface
    input             CF_cfgb_awvalid,        // Write Address Valid
    output            BC_cfgb_awready,        // Write Address Port Ready
    input      [23:0] CF_cfgb_awaddr,         // Write Address
    input             CF_cfgb_wvalid,         // Write Data Valid
    output            BC_cfgb_wready,         // Write Data Port Ready
    input      [31:0] CF_cfgb_wdata,          // Write Data
    input      [3:0]  CF_cfgb_wstrb,          // Write Data Byte Enables
    output            BC_cfgb_bvalid,         // Write Response Valid
    input             CF_cfgb_bready,         // Write Response Fabric Ready
    input             CF_cfgb_arvalid,        // Read Address Valid
    output            BC_cfgb_arready,        // Read Address Port Ready
    input      [23:0] CF_cfgb_araddr,         // Read Address
    output            BC_cfgb_rvalid,         // Read Response Valid
    input             CF_cfgb_rready,         // Read Response Fabric Ready
    output     [31:0] BC_cfgb_rdata           // Read Data
    // }}} End Port Declarations -----------
  );

  // {{{ Wire Declarations -----------------
  wire                CCA_sync_cfg_rst;       // cfg_rst sync'ed to phy_clk
  wire         [23:0] CCA_cfg_waddr;          // Write Address
  wire         [31:0] CCA_cfg_wdata;          // Write Data
  wire         [3:0]  CCA_cfg_wstrb;          // Write Data Byte Enables
  wire                CCA_sync_we;            // Synchronized write enable
  wire         [23:0] CCA_cfg_raddr;          // Read Address
  wire                CCA_sync_re;            // Synchronized Read Enable
  wire         [31:0] BCR_core_rdata;         // Read Data
  // }}} End Wire Declarations -------------


  // {{{ cfg_axi Inst ----------------------
  // Instantiate the generic cfg interface, which contains the clock domain
  // crossing from cfg_clk to phy_clk, as well as the
  // AXI-Lite interface to the CFG Fabric
  srio_gen2_v4_1_16_cfg_axi
    #(
      .TCQ                       (TCQ))
    buf_cfg_axi_inst
     (.core_clk                  (phy_clk),
      .cfg_clk                   (cfg_clk),
      .cfg_rst                   (cfg_rst),
      .CF_awvalid                (CF_cfgb_awvalid),
      .CCA_awready               (BC_cfgb_awready),
      .CF_awaddr                 (CF_cfgb_awaddr),
      .CF_wvalid                 (CF_cfgb_wvalid),
      .CCA_wready                (BC_cfgb_wready),
      .CF_wdata                  (CF_cfgb_wdata),
      .CF_wstrb                  (CF_cfgb_wstrb),
      .CCA_bvalid                (BC_cfgb_bvalid),
      .CF_bready                 (CF_cfgb_bready),
      .CF_arvalid                (CF_cfgb_arvalid),
      .CCA_arready               (BC_cfgb_arready),
      .CF_araddr                 (CF_cfgb_araddr),
      .CCA_rvalid                (BC_cfgb_rvalid),
      .CF_rready                 (CF_cfgb_rready),
      .CCA_rdata                 (BC_cfgb_rdata),
      .CCA_sync_cfg_rst          (CCA_sync_cfg_rst),
      .CCA_cfg_waddr             (CCA_cfg_waddr),
      .CCA_cfg_wdata             (CCA_cfg_wdata),
      .CCA_cfg_wstrb             (CCA_cfg_wstrb),
      .CCA_sync_we               (CCA_sync_we),
      .CCA_cfg_raddr             (CCA_cfg_raddr),
      .CCA_sync_re               (CCA_sync_re),
      .CC_core_rdata             (BCR_core_rdata));
  // }}} End cfg_axi Inst ------------------

  // {{{ buf_cfg_reg Inst ------------------
  // Instantiate the BUF CFG register bank, containing all the CSRs for the Buffer
  srio_gen2_v4_1_16_buf_cfg_reg
    #(
      .TCQ                       (TCQ),
      .TX_DEPTH                  (TX_DEPTH),
      .RX_DEPTH                  (RX_DEPTH),
      .RX_FC_ONLY                (RX_FC_ONLY),
      .UNIFIED_CLK               (UNIFIED_CLK),
      .REQ_REORDER               (REQ_REORDER),
      .WM0                       (WM0),
      .WM1                       (WM1),
      .WM2                       (WM2),
      .IDLE2                     (IDLE2))
  buf_cfg_reg_inst
    (
      .phy_clk                   (phy_clk),
      .buf_phy_rst               (buf_phy_rst),
      .CCA_sync_cfg_rst          (CCA_sync_cfg_rst),
      .BT_tx_flow_control        (BT_tx_flow_control),
      .PP_idle2_selected         (PP_idle2_selected),
      .BCR_watermark0            (BC_watermark0),
      .BCR_watermark1            (BC_watermark1),
      .BCR_watermark2            (BC_watermark2),
      .BCR_force_rx_flow         (BC_force_rx_flow),
      .CCA_cfg_waddr             (CCA_cfg_waddr),
      .CCA_cfg_wdata             (CCA_cfg_wdata),
      .CCA_cfg_wstrb             (CCA_cfg_wstrb),
      .CCA_sync_we               (CCA_sync_we),
      .CCA_cfg_raddr             (CCA_cfg_raddr),
      .CCA_sync_re               (CCA_sync_re),
      .BCR_core_rdata            (BCR_core_rdata));
  // }}} End buf_cfg_reg Inst --------------

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/buf/buf_cfg/srio_gen2_v4_1_16_buf_cfg_reg.v#1 $
//----------------------------------------------------------------------
//
// BUF_CFG_REG
// Description:
// This module contains the configuration registers for the Buffer.
//
// For writes, it takes a write enable, address, data and strobe (byte
// enables) from the cfg_axi module, decodes the address, and updates
// applicable registers. For reads, it takes an address and read enable,
// and returns the read data from the corresponding CSR. It also has a
// buffer core interface for transfer of control and status information.
//
// No clock relationship between the cfg_clk and the phy_clk is assumed.
//
// Hierarchy:
// BUF_TOP
//    |______BUF_CFG_TOP
//              |______CFG_AXI (in hdl/common/)
//              |______BUF_CFG_REG <-- this module
// ---------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)

module srio_gen2_v4_1_16_buf_cfg_reg
  #(
    parameter TCQ         = 100,
    parameter TX_DEPTH    = 32,   // TX buffer depth {8, 16, 32}
    parameter RX_DEPTH    = 32,   // RX buffer depth {8, 16, 32}
    parameter RX_FC_ONLY  = 0,    // RX Flow Control Only {0, 1}
    parameter UNIFIED_CLK = 0,    // phy_clk = log_clk {0, 1}
    parameter REQ_REORDER = 1,    // Request reordering enabled {0, 1}
    parameter WM0         = 3,    // Watermark 0 reset value {WM0 < 64}
    parameter WM1         = 2,    // Watermark 1 reset value {WM0 > WM1 > WM2}
    parameter WM2         = 1,    // Watermark 2 reset value {WM2 > 0}
    parameter IDLE2       = 0)    // IDLE2 sequence support
  (
    // {{{ Port Declarations ---------------
    // System Signals
    input             phy_clk,                        // PHY interface clock
    input             buf_phy_rst,                    // Reset for PHY clock Domain
    input             CCA_sync_cfg_rst,               // cfg_rst sync'ed to phy_clk

    // Buffer Interface 
    // Initialize signals going to buffer that are reset on CCA_sync_cfg_rst to avoid sim X's
    input             BT_tx_flow_control,             // TX Flow Control Mode
    input             PP_idle2_selected,              // OPLM has trained to use IDLE2 sequence
    output reg [5:0]  BCR_watermark0 = WM0,           // Watermark 0
    output reg [5:0]  BCR_watermark1 = WM1,           // Watermark 1
    output reg [5:0]  BCR_watermark2 = WM2,           // Watermark 2
    output reg        BCR_force_rx_flow = RX_FC_ONLY, // Force the Buffer into RX Flow Control mode

    // Generic Configuration Interface
    input      [23:0] CCA_cfg_waddr,                  // Write Address
    input      [31:0] CCA_cfg_wdata,                  // Write Data
    input      [3:0]  CCA_cfg_wstrb,                  // Write Data Byte Enables
    input             CCA_sync_we,                    // Synchronized write enable
    input      [23:0] CCA_cfg_raddr,                  // Read Address
    input             CCA_sync_re,                    // Synchronized Read Enable
    output reg [31:0] BCR_core_rdata                  // Read Data
    // }}} End Port Declarations -----------
  );

  // {{{ Localparams -----------------------
  localparam [5:0]  WM0_MAX   = 6'd29;        // Max value for WM0 when IDLE1 sequence in use
  localparam [5:0]  WM1_MAX   = 6'd28;        // Max value for WM1 when IDLE1 sequence in use
  localparam [5:0]  WM2_MAX   = 6'd27;        // Max value for WM2 when IDLE1 sequence in use
  
  // Parameters for CSR offsets
  // It is assumed that the MSB of the address for received reads and writes matches the buffer config offset
  localparam [15:0] BUF_000   = 16'h0000;   // Watermarks CSR
  localparam [15:0] BUF_004   = 16'h0004;   // Buffer Control CSR
  // }}} End Localparams -------------------

  // {{{ Wire Declarations -----------------
  reg           tx_flow_control;              // registered version of BT_tx_flow_control for fanout control
  wire  [31:0]  csr_buf_000, csr_buf_004;     // wires representing each CSR for ease of use in simulation
  reg   [5:0]   buf_000_wm0;                  // Written watermark 0 value
  reg   [5:0]   buf_000_wm1;                  // Written watermark 1 value
  reg   [5:0]   buf_000_wm2;                  // Written watermark 2 value
  // }}} End Wire Declarations -------------
  
  // {{{ Core Fanout Control ---------------
  always @(posedge phy_clk) begin
    // Unnecessary to have reset value since it's assigned from inputs
    // on every cycle 
    tx_flow_control   <= #TCQ BT_tx_flow_control;
  end
  // }}} End Core Fanout Control -----------
  
  
  // {{{ Writable Register Bank ------------
  // A shadow register is kept for writable registers so that read and write 
  // functionality can be fully separated.
  // ----- Port Link Timeout CSR writable register(s) ----- //
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      buf_000_wm2           <= #TCQ WM2;
      buf_000_wm1           <= #TCQ WM1;
      buf_000_wm0           <= #TCQ WM0;
    end else if (CCA_sync_we && (CCA_cfg_waddr[15:0] == BUF_000)) begin
      if (IDLE2 == 1) begin
        if (CCA_cfg_wstrb[2])
          buf_000_wm2       <= #TCQ CCA_cfg_wdata[21:16];
        if (CCA_cfg_wstrb[1])
          buf_000_wm1       <= #TCQ CCA_cfg_wdata[13:8];
        if (CCA_cfg_wstrb[0])
          buf_000_wm0       <= #TCQ CCA_cfg_wdata[5:0];
      end else begin
        if (CCA_cfg_wstrb[2])
          buf_000_wm2       <= #TCQ {1'b0, CCA_cfg_wdata[20:16]};
        if (CCA_cfg_wstrb[1])
          buf_000_wm1       <= #TCQ {1'b0, CCA_cfg_wdata[12:8]};
        if (CCA_cfg_wstrb[0])
          buf_000_wm0       <= #TCQ {1'b0, CCA_cfg_wdata[4:0]};
      end
    end
  end
  
  //*COVERAGE*
  //(cp_wm0): Cover various values written for WM0

  //*COVERAGE*
  //(cp_wm1): Cover various values written for WM1

  //*COVERAGE*
  //(cp_wm2): Cover various values written for WM2
    
  // Create watermark outputs
  // If IDLE2 is not supported, the watermarks are 5 bits and the user is expected to write valid values.
  // If IDLE2 is supported, the watermarks are 6 bits. If the OPLM trains to use IDLE1, we'll limit the 
  // watermarks to their practical maximums to avoid the possibility of locking up the TX buffer. The CSR
  // will still return the last written value when read.
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      BCR_watermark2        <= #TCQ WM2;
      BCR_watermark1        <= #TCQ WM1;
      BCR_watermark0        <= #TCQ WM0;
    end else if (IDLE2 == 0) begin
      BCR_watermark2        <= #TCQ buf_000_wm2;
      BCR_watermark1        <= #TCQ buf_000_wm1;
      BCR_watermark0        <= #TCQ buf_000_wm0;
    end else if (PP_idle2_selected) begin
      BCR_watermark2        <= #TCQ buf_000_wm2;
      BCR_watermark1        <= #TCQ buf_000_wm1;
      BCR_watermark0        <= #TCQ buf_000_wm0;
    // If IDLE2 is supported but the OPLM has trained to use IDLE1 sequence, limit the watermark values to the buffer
    end else begin // Should only be hit if !CCA_sync_cfg_rst && !PP_idle2_selected && (IDLE2 == 1)
      BCR_watermark2        <= #TCQ ((buf_000_wm2 > WM2_MAX) ? WM2_MAX : buf_000_wm2);
      BCR_watermark1        <= #TCQ ((buf_000_wm1 > WM1_MAX) ? WM1_MAX : buf_000_wm1);
      BCR_watermark0        <= #TCQ ((buf_000_wm0 > WM0_MAX) ? WM0_MAX : buf_000_wm0);
    end
  end

  // ----- Port Response Timeout CSR writable register(s) ----- //
  always @(posedge phy_clk) begin
    if (CCA_sync_cfg_rst) begin
      BCR_force_rx_flow     <= #TCQ RX_FC_ONLY;
    end else if (RX_FC_ONLY == 1) begin
      BCR_force_rx_flow     <= #TCQ RX_FC_ONLY;
    end else if (CCA_sync_we && (CCA_cfg_waddr[15:0] == BUF_004)) begin
      if (CCA_cfg_wstrb[1])
        BCR_force_rx_flow   <= #TCQ CCA_cfg_wdata[15];
    end
  end

  //*COVERAGE*
  //(cp_force_rx_flow): Enumerate the value written for force_rx_flow
  
  // }}} End Writable Register Bank ---------

  
  
  // {{{ Read Data Assembly ----------------
  // Form read data based on address
  // Bit ordering mirrors RapidIO Spec (e.g. spec bit 0 -> phy_cfg bit 31)
  
  // Create wires for each CSR for easy simulation viewing.
  
  // ------------------- Buffer Configuration Registers ---------------------------
                                                    // core  (spec)   Description
                                                    // ----------------------------
  // Watermarks CSR
  assign csr_buf_000 =  {10'b0,                     // 31:22  (0:9)   Reserved
                         buf_000_wm2,               // 21:16  (10:15) Watermark 2
                         2'b0,                      // 15:14  (16:17) Reserved
                         buf_000_wm1,               // 13:8   (18:23) Watermark 1
                         2'b0,                      // 7:6    (24:25) Reserved
                         buf_000_wm0};              // 5:0    (26:31) Watermark 0
                         
  // Buffer Control CSR
  assign csr_buf_004 =  {(RX_FC_ONLY == 1),         // 31     (0)     RX Flow Control Only
                         (UNIFIED_CLK == 1),        // 30     (1)     Unified Clock
                         tx_flow_control,           // 29     (2)     TX Flow Control
                         (REQ_REORDER == 1),        // 28     (3)     Request Reorder Support
                         4'b0,                      // 27:24  (4:7)   Reserved
                         TX_DEPTH[7:0],             // 23:16  (8:15)  TX Size
                         BCR_force_rx_flow,         // 15     (16)    Force RX Flow Control
                         7'b0,                      // 14:8   (17:23) Reserved
                         RX_DEPTH[7:0]};            // 7:0    (24:31) RX Size

  //*COVERAGE*
  //(cp_buf_000_3_rd_b4_wr): Cover that buf_000 byte 3 was read before it was written
  //(cp_buf_000_2_rd_b4_wr): Cover that buf_000 byte 2 was read before it was written
  //(cp_buf_000_1_rd_b4_wr): Cover that buf_000 byte 1 was read before it was written
  //(cp_buf_000_0_rd_b4_wr): Cover that buf_000 byte 0 was read before it was written
  //(cp_buf_000_3_rd_aftr_wr): Cover that buf_000 byte 3 was read after it was written
  //(cp_buf_000_2_rd_aftr_wr): Cover that buf_000 byte 2 was read after it was written
  //(cp_buf_000_1_rd_aftr_wr): Cover that buf_000 byte 1 was read after it was written
  //(cp_buf_000_0_rd_aftr_wr): Cover that buf_000 byte 0 was read after it was written
  //(cp_buf_000_2_rst_val_chk): Cover that WM2 is non-default and buf_000 byte 2 was rd_b4_wr
  //(cp_buf_000_1_rst_val_chk): Cover that WM1 is non-default and buf_000 byte 1 was rd_b4_wr
  //(cp_buf_000_0_rst_val_chk): Cover that WM0 is non-default and buf_000 byte 0 was rd_b4_wr
  //(cp_buf_004_3_rd_b4_wr): Cover that buf_004 byte 3 was read before it was written
  //(cp_buf_004_2_rd_b4_wr): Cover that buf_004 byte 2 was read before it was written
  //(cp_buf_004_1_rd_b4_wr): Cover that buf_004 byte 1 was read before it was written
  //(cp_buf_004_0_rd_b4_wr): Cover that buf_004 byte 0 was read before it was written
  //(cp_buf_004_3_rd_aftr_wr): Cover that buf_004 byte 3 was read after it was written
  //(cp_buf_004_2_rd_aftr_wr): Cover that buf_004 byte 2 was read after it was written
  //(cp_buf_004_1_rd_aftr_wr): Cover that buf_004 byte 1 was read after it was written
  //(cp_buf_004_0_rd_aftr_wr): Cover that buf_004 byte 0 was read after it was written
  //(cp_buf_004_bit31_rst_val_chk): Cover that RX_FC_ONLY is non-default and buf_004 bit 31 was rd_b4_wr
  //(cp_buf_004_bit30_rst_val_chk): Cover that UNIFIED_CLK is non-default and buf_004 bit 30 was rd_b4_wr
  //(cp_buf_004_bit28_rst_val_chk): Cover that REQ_REORDER is non-default and buf_004 bit 28 was rd_b4_wr
  //(cp_buf_004_2_rst_val_chk): Cover that TX_DEPTH is non-default and buf_004 byte 2 was rd_b4_wr
  //(cp_buf_004_0_rst_val_chk): Cover that RX_DEPTH is non-default and buf_004 byte 2 was rd_b4_wr

  // Register read data when address is safe
  // No reset needed since data is not sampled until valid
  always @(posedge phy_clk) begin
    if (CCA_sync_re) begin
      case (CCA_cfg_raddr[15:0])
        BUF_000    : BCR_core_rdata <= #TCQ csr_buf_000;
        BUF_004    : BCR_core_rdata <= #TCQ csr_buf_004;
        // Return data of all 0's if read to unimplemented space
        default    : BCR_core_rdata <= #TCQ 32'b0;      
      endcase
    end
  end

  // }}} End Read Data Assembly ------------
  

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/buf/srio_gen2_v4_1_16_buf_rx_bram_bank.v#1 $
//
// BUF_RX_BRAM_BANK
// Description:
// This module instantiates a family-specific memory module. It calls
// BLK_MEM_GEN from Coregen
//
// Hierarchy:
// BUF_TOP
//  |______BUF_TX
//  |____________BUF_TX_SYNC_UNIT
//  |____________BUF_TX_BRAM_BANK
//  |______BUF_RX
//  |____________BUF_RX_ASYNC_PASSAGE
//  |____________BUF_RX_BRAM_BANK <-- this module
//----------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)


module srio_gen2_v4_1_16_buf_rx_bram_bank
  #(
    parameter TCQ           = 100,
    parameter UNIFIED_CLK   = 0,                 // {0, 1}
    parameter C_FAMILY      = "virtex6",         // {virtex5, virtex6, virtex7, spartan6, spartan7}
    parameter C_ADDR_LEN    = 11)                // {9, 10, 11}
   (
   // {{{ port declarations -----------------
    input                   phy_clk,             // Physical Layer clock
    input                   log_clk,             // Logical Layer clock
    input                   buf_phy_rst_q,       // Synchronous Phy Layer reset
    input                   buf_log_rst_q,       // Synchronous Log Layer reset
    // in from Physical clock
    input  [C_ADDR_LEN-1:0] BR_phy_bram_waddr,   // Write address for memory
    input                   BR_phy_bram_we,      // Write enable
    input  [63:0]           PR_phy_tdata_q,      // Data In
    input  [1:0]            PR_phy_tuser_q,      // User Field
    input  [2:0]            PR_phy_tkeep_q,      // Remainder
    input                   PR_phy_tlast_q,      // End of Frame
    // in/out to Logical clock
    input  [C_ADDR_LEN-1:0] BR_log_bram_raddr,   // Read address for memory
    input                   BR_log_bram_rd,      // Read enable
    output [63:0]           BRB_log_bram_tdata,  // Data Out
    output [1:0]            BRB_log_bram_tuser,  // Critical Request Flow
    output [2:0]            BRB_log_bram_tkeep,  // Remainder
    output                  BRB_log_bram_tlast   // End of Frame
   // }}} ---------------------------------
   );


  // {{{ local parameters ------------------
  localparam C_MEM_DEPTH = 1 << C_ADDR_LEN;
  // }}} ---------------------------------

  // {{{ wire declarations -----------------
  wire [69:0] bram_data_in  = {PR_phy_tlast_q, PR_phy_tkeep_q, PR_phy_tuser_q, PR_phy_tdata_q};
  wire [69:0] bram_data_out;

  assign {BRB_log_bram_tlast, BRB_log_bram_tkeep, BRB_log_bram_tuser, BRB_log_bram_tdata}  = bram_data_out;

//  assign BRB_log_bram_tlast  = bram_data_out[69];
//  assign BRB_log_bram_tkeep  = bram_data_out[68:66];
//  assign BRB_log_bram_tuser  = bram_data_out[65:64];
//  assign BRB_log_bram_tdata  = bram_data_out[63:0];
  // }}} ---------------------------------

  // {{{ Block memory Instantiation --------
  blk_mem_gen_v8_4_4                                       // blk_mem_gen_v8_0 values 
   #(
     .C_ADDRA_WIDTH               (C_ADDR_LEN),          // (C_ADDR_LEN),
     .C_ADDRB_WIDTH               (C_ADDR_LEN),          // (C_ADDR_LEN),
     .C_ALGORITHM                 (1),                   // (1),
     .C_AXI_ID_WIDTH              (4),                   // (4),
     .C_AXI_SLAVE_TYPE            (4), //(0),            // (4),
     .C_AXI_TYPE                  (4), //(1),            // (4),
     .C_BYTE_SIZE                 (9),                   // (9),
     .C_COMMON_CLK                (UNIFIED_CLK),         // (UNIFIED_CLK),
     .C_DEFAULT_DATA              ("0"),                 // ("0"),
     .C_DISABLE_WARN_BHV_COLL     (0),                   // (0),
     .C_DISABLE_WARN_BHV_RANGE    (1),                   // (1),
     .C_ELABORATION_DIR           ("./"),                // (""),
     .C_ENABLE_32BIT_ADDRESS      (0),                   // (0),
     .C_FAMILY                    (C_FAMILY),            // (C_FAMILY),
     .C_HAS_AXI_ID                (0),                   // (0),
     .C_HAS_ENA                   (1),                   // (1),
     .C_HAS_ENB                   (1),                   // (1),
     .C_HAS_INJECTERR             (0),                   // (0),
     .C_HAS_MEM_OUTPUT_REGS_A     (0),                   // (0),
     .C_HAS_MEM_OUTPUT_REGS_B     (1),                   // (1),
     .C_HAS_MUX_OUTPUT_REGS_A     (0),                   // (0),
     .C_HAS_MUX_OUTPUT_REGS_B     (0),                   // (0),
     .C_HAS_REGCEA                (0),                   // (0),
     .C_HAS_REGCEB                (0),                   // (0),
     .C_HAS_RSTA                  (0),//(1),             // (0),
     .C_HAS_RSTB                  (1),                   // (1),
     .C_HAS_SOFTECC_INPUT_REGS_A  (0),                   // (0),
     .C_HAS_SOFTECC_OUTPUT_REGS_B (0),                   // (0),
     .C_INIT_FILE_NAME            ("no_coe_file_loaded"),// ("no_coe_file_loaded"),
     .C_INITA_VAL                 ("0"),                 // ("0"),
     .C_INITB_VAL                 ("0"),                 // ("0"),
     .C_INTERFACE_TYPE            (0),                   // (0),
     .C_LOAD_INIT_FILE            (0),                   // (0),
     .C_MEM_TYPE                  (1),                   // (1),
     .C_MUX_PIPELINE_STAGES       (0),                   // (0),
     .C_PRIM_TYPE                 (1),                   // (1),
     .C_READ_DEPTH_A              (C_MEM_DEPTH),         // (C_MEM_DEPTH),
     .C_READ_DEPTH_B              (C_MEM_DEPTH),         // (C_MEM_DEPTH),
     .C_READ_WIDTH_A              (70),                  // (70),
     .C_READ_WIDTH_B              (70),                  // (70),
     .C_RST_PRIORITY_A            ("CE"),                // ("CE"),
     .C_RST_PRIORITY_B            ("CE"),                // ("CE"),
     //.C_RST_TYPE                  ("SYNC"),              // ("SYNC"),// removed in v8_2 instance
     .C_RSTRAM_A                  (0),                   // (0),
     .C_RSTRAM_B                  (0),                   // (0),
     .C_SIM_COLLISION_CHECK       ("NONE"),              // ("NONE"),
     .C_USE_BYTE_WEA              (0),                   // (0),
     .C_USE_BYTE_WEB              (0),                   // (0),
     .C_USE_DEFAULT_DATA          (0),                   // (0),
     .C_USE_ECC                   (0),                   // (0),
     .C_USE_SOFTECC               (0),                   // (0),
     .C_WEA_WIDTH                 (1),                   // (1),
     .C_WEB_WIDTH                 (1),                   // (1),
     .C_WRITE_DEPTH_A             (C_MEM_DEPTH),         // (C_MEM_DEPTH),
     .C_WRITE_DEPTH_B             (C_MEM_DEPTH),         // (C_MEM_DEPTH),
     .C_WRITE_MODE_A              ("WRITE_FIRST"),       // ("WRITE_FIRST"),
     .C_WRITE_MODE_B              ("WRITE_FIRST"),       // ("WRITE_FIRST"),
     .C_WRITE_WIDTH_A             (70),                  // (70),
     .C_WRITE_WIDTH_B             (70),                  // (70),
     .C_XDEVICEFAMILY             (C_FAMILY),            // (C_FAMILY))

     // newly added parameters for the Diablo/US updates, leave default // 1/13/2015
     .C_USE_URAM                    (0),
     .C_EN_SAFETY_CKT               (0),
     .C_EN_DEEPSLEEP_PIN	    (0),
     .C_EN_SHUTDOWN_PIN	            (0),
     .C_EN_RDADDRA_CHG	            (0),
     .C_EN_RDADDRB_CHG	            (0)

     //_____________Below are newly added with blk_mem_gen_v8_2 version
     //_____________as per block mem gen owner, can be left at default or
     //_____________not included in the instance
     // .C_USE_BRAM_BLOCK		(0),
     // .C_CTRL_ECC_ALGO		("NONE"),
     // .C_INIT_FILE		("blk_mem_gen_0.mem"),
     // .C_EN_ECC_PIPE		(0),
     // .C_EN_SLEEP_PIN		(0),
     // .C_COUNT_36K_BRAM		("0"),
     // .C_COUNT_18K_BRAM		("1"),
     // .C_EST_POWER_SUMMARY	("Estimated Power for IP     :     3.0361 mW")
     )            
   blk_mem_inst
    (.clka                        (phy_clk),
     .dina                        (bram_data_in),
     .addra                       (BR_phy_bram_waddr),
     .ena                         (1'b1),
     .regcea                      (1'b0),
     .wea                         (BR_phy_bram_we),
     .rsta                        (buf_phy_rst_q),
     .douta                       (),
     .clkb                        (log_clk),
     .dinb                        (70'h0),
     .addrb                       (BR_log_bram_raddr),
     .enb                         (BR_log_bram_rd),
     .regceb                      (1'b0),
     .web                         (1'b0),
     .rstb                        (buf_log_rst_q),
     .doutb                       (bram_data_out),
     .sbiterr                     (),
     .dbiterr                     (),
     .injectsbiterr               (),
     .injectdbiterr               (),
     .rdaddrecc                   (),

   // dont touch ports, new addition with default drive, // 1/13/2015
     .deepsleep                   (1'b0),
     .shutdown                    (1'b0),

     .s_aclk                      (),
     .s_aresetn                   (),
     .s_axi_awid                  (),
     .s_axi_awaddr                (),
     .s_axi_awlen                 (),
     .s_axi_awsize                (),
     .s_axi_awburst               (),
     .s_axi_awvalid               (),
     .s_axi_awready               (),
     .s_axi_wdata                 (),
     .s_axi_wstrb                 (),
     .s_axi_wlast                 (),
     .s_axi_wvalid                (),
     .s_axi_wready                (),
     .s_axi_bid                   (),
     .s_axi_bresp                 (),
     .s_axi_bvalid                (),
     .s_axi_bready                (),
     .s_axi_arid                  (),
     .s_axi_araddr                (),
     .s_axi_arlen                 (),
     .s_axi_arsize                (),
     .s_axi_arburst               (),
     .s_axi_arvalid               (),
     .s_axi_arready               (),
     .s_axi_rid                   (),
     .s_axi_rdata                 (),
     .s_axi_rresp                 (),
     .s_axi_rlast                 (),
     .s_axi_rvalid                (),
     .s_axi_rready                (),
     .s_axi_injectsbiterr         (),
     .s_axi_injectdbiterr         (),
     .s_axi_sbiterr               (),
     .s_axi_dbiterr               (),
     .s_axi_rdaddrecc             (),
     .sleep                       (1'b0),
     .eccpipece                   (1'b0)
    );
  // }}} ---------------------------------

endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/buf/srio_gen2_v4_1_16_buf_rx.v#1 $
//
// BUF_RX
// Description:
// This module is the RX path of the BUFFER. It is responsible for the 
// following:
// 1. Receiving Data from the Physical Layer
// 2. Storing and packets until delivery to the Logical Layer
//   
// Hierarchy:
// BUF_TOP
//  |______BUF_TX
//  |____________BUF_TX_SYNC_UNIT
//  |____________BUF_TX_BRAM_BANK
//  |______BUF_RX <-- this module
//  |____________BUF_RX_ASYNC_PASSAGE
//  |____________BUF_RX_BRAM_BANK
//----------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)

module srio_gen2_v4_1_16_buf_rx
  #(
    parameter TCQ           = 100,
    parameter MODE_XG       = 5,           // {1, 2, 3, 5, 6}
    parameter HW_ARCH       = 2,           // {0 -8} indication of architecture
    parameter RX_DEPTH      = 32,          // {8, 16, 32}
    parameter UNIFIED_CLK   = 0,           // {0, 1}
    parameter EVAL          = 1)           // {0, 1}
   (
    // {{{ port declarations ---------------
    // clocks and resets
    input             log_clk,             // Freerunning Logical Layer clock
    input             phy_clk,             // Freerunning Physical Layer clock
    input             buf_log_rst,         // Synchronous Logical Layer reset
    input             buf_phy_rst,         // Synchronous Physical Layer reset

    // LOG RX Interface
    output reg        BR_bufr_tvalid,      // Valid Packet Beat
    input             LE_bufr_tready,      // Packet Beat Accepted
    output reg [63:0] BR_bufr_tdata,       // Packet Data
    output reg  [7:0] BR_bufr_tkeep,       // Valid bytes in this beat, only valid on last
    output reg        BR_bufr_tlast,       // Last Beat
    output reg  [7:0] BR_bufr_tuser,       // {4'h0, SOP, VC, CRF, 1'b0} AXI Compliance Pad

    // PHY RX Interface
    input             PR_phyr_tvalid,      // Valid Data Indicator
    output reg        BR_phyr_tready,      // Destination Ready
    input      [63:0] PR_phyr_tdata,       // Packet Data
    input       [7:0] PR_phyr_tkeep,       // Byte Enable for Data, only valid on last
    input             PR_phyr_tlast,       // Last DW of Packet Data
    input       [7:0] PR_phyr_tuser,       // {5'h00, VC, CRF, src_dsc} AXI Compliance Pad
    output reg  [5:0] BR_phy_buf_stat      // Buffer Status from the RX Buffer
    // }}} ---------------------------------
   );


  // {{{ local parameters ----------------

  // Since the RX buffer doesn't segment BRAM the same way as TX,
  // RX_DEPTH does not indicate a true number of packets that can be stored
  // for a given configuration. It is being kept to match the notation of
  // of the TX buffer. Instead, a value of 8 occupies 1 BRAM, 16 occupies 2,
  // 32 occupies 4. Each value of RX_DEPTH can store at least that many max-sized
  // packets (and likely many more).
  localparam       C_TAG_LEN   = RX_DEPTH ==  8 ? 3 :
                                 RX_DEPTH == 16 ? 4 :
                                 RX_DEPTH == 32 ? 5 :
                                                  1; // undefined
  localparam [2:0] C_MAX_INDEX_LEN = 6;
  localparam [3:0] C_ADDR_LEN      = C_TAG_LEN + C_MAX_INDEX_LEN;

  localparam       C_FAMILY    = HW_ARCH == 0 ? "virtex5"  :
                                 HW_ARCH == 1 ? "virtex5"  :
                                 HW_ARCH == 2 ? "virtex6"  :
                                 HW_ARCH == 3 ? "virtex6"  :
                                 HW_ARCH == 4 ? "spartan6" :
                                 HW_ARCH == 5 ? "artix7"   :
                                 HW_ARCH == 6 ? "kintex7"  :
                                 HW_ARCH == 7 ? "virtex7"  :
                                 HW_ARCH == 8 ? "virtex7"  :
                                 HW_ARCH == 9 ? "zynq"  :
                                 HW_ARCH == 10 ? "ultrascale"  :
                                 HW_ARCH == 11 ? "ultrascale"  :
                                 HW_ARCH == 12 ? "ultrascale"  :
                                 HW_ARCH == 13 ? "ultrascale"  :
                                 HW_ARCH == 14 ? "ultrascale"  :
                                                "undefined";

// added below macro to fix the CR# 735137
// synthesis translate_off 
  initial begin
    if (C_TAG_LEN == 1) begin
      $display("ERROR: RX_DEPTH holds an unexpected value in buf_rx");
      $finish;
    end
    if (C_FAMILY == "undefined") begin
      $display("ERROR: HW_ARCH holds an unexpected value in buf_rx");
      $finish;
    end
  end
  // }}} ---------------------------------
// synthesis translate_on

  // {{{ wire declarations ---------------
  // Prefix notation:
  // phy = phy clock domain
  // log = log clock domain
  // bufr = AXI LOG - BUF interface
  // phyr = AXI PHY - BUF interface
  // pr/PR = Physical Layer Receive (only used on ports)
  // br/BR = Buffer Layer Receive (only used on ports)
  // brp = Async Passage within Receive Buffer (only used on ports)
  // brb = BRAM Bank within Receive Buffer (only used on ports)

  // resets
  reg                    buf_phy_rst_q = 1;       // registered physical layer reset
  reg                    buf_log_rst_q = 1;       // registered logical layer reset

  // PHY clock domain signals
  reg                    pr_phyr_tlast_q;         // registered only when valid
  reg  [63:0]            pr_phyr_tdata_q;         // registered only when valid
  reg   [2:0]            pr_phyr_tkeep_q;         // reduced version of the actual strobe
  reg   [1:0]            pr_phyr_tuser_q;         // only stores VC and CRF bits
  reg                    pr_phyr_src_dsc_q;       // registered source discontinue
  wire                   phy_phase_valid;         // indicates a valid data beat within a packet
  wire                   complete_packet_written; // a packet has been stored succesfully w/o discontinue
  wire [C_ADDR_LEN-1:0]  brp_phy_bram_raddr;      // read address converted to the phy domain

  // BRAM Bank signals
  reg                    br_phy_bram_we;          // buffer write enable
  reg  [C_ADDR_LEN-1:0]  br_phy_bram_waddr;       // buffer write address

  wire                   br_log_bram_rd;          // buffer read enable
  reg  [C_ADDR_LEN-1:0]  br_log_bram_raddr;       // buffer read address
  wire [63:0]            brb_log_bram_tdata;      // buffered data output
  wire [1:0]             brb_log_bram_tuser;      // buffered data output
  wire [2:0]             brb_log_bram_tkeep;      // buffered data output
  wire                   brb_log_bram_tlast;      // buffered data output

  // LOG clock domain signals
  wire [C_ADDR_LEN-1:0]  brp_log_starting_waddr;  // log domain number of packets written into buffer 
  reg                    log_set_empty_condition; // asserts when it appears that the buffer goes empty
  wire                   log_set_empty;           // set buffer empty
  wire                   log_clr_empty;           // clear buffer empty
  wire                   log_pipeline_vacancy;    // when asserted, there is a free location in the pipe
  reg  [1:0]             log_pipeline_count;      // counts the number of data beats in the pipeline
  reg  [1:0]             br_bufr_tvalid_d;        // coincides with internal pipeline stages
  reg                    buf_tstart;              // This is the REAL SOP, embedded into TUSER
  reg                    buf_log_sof_out;         // This is the timeout circuit output
  wire                   buf_log_sof_out_d;       // This is the timeout circuit output
  reg                    log_buffer_empty;        // buffer empty indication
  reg                    br_bufr_tvalid_q;        // registered version of tvalid

  // }}} ---------------------------------


  // {{{ Reset Structure -----------------

  // by rule, we must register the resets before we use them. This is not a
  // synchronizing circuit but rather a method to reduce fanout on the resets.
  //always @(posedge phy_clk or posedge buf_phy_rst) begin
  always @(posedge phy_clk) begin
    if (buf_phy_rst)
      buf_phy_rst_q <= #TCQ 1'b1;
    else
      buf_phy_rst_q <= #TCQ 1'b0;
  end
  //always @(posedge log_clk or posedge buf_log_rst) begin
  always @(posedge log_clk ) begin
    if (buf_log_rst)
      buf_log_rst_q <= #TCQ 1'b1;
    else
      buf_log_rst_q <= #TCQ 1'b0;
  end


    // *- ASSERTION (BR_reset_behavior)
    // buf_log_rst and buf_phy_rst must overlap when driven high.

  // }}} ---------------------------------


  // {{{ PHY Interface -------------------
  assign phy_phase_valid = PR_phyr_tvalid && BR_phyr_tready;

  // capture data only on valid data beats. Use resets on the control signals. Data doesn't need reset.
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      pr_phyr_tlast_q   <= #TCQ 1'b0;
      pr_phyr_src_dsc_q <= #TCQ 1'b0;
    end else if (phy_phase_valid) begin
      pr_phyr_tlast_q   <= #TCQ PR_phyr_tlast;
      pr_phyr_src_dsc_q <= #TCQ PR_phyr_tuser[0];
    end
  end
  always @(posedge phy_clk) begin
    if (phy_phase_valid) begin
      pr_phyr_tdata_q   <= #TCQ PR_phyr_tdata;
      pr_phyr_tuser_q   <= #TCQ PR_phyr_tuser[2:1];
    end
  end

  // 3 bit encoding for tkeep. There are only four valid remainder combinations when tlast is asserted.
  // Just grab every other value, which is enough to reconstruct the strobe on the other end.
  // NOTE: when reconstructing, it is expected that strobe be FF when in a packet other than the last beat.
  // There is an assertion to make sure this happenen in the IF bind. Otherwise, the reconstruction on the
  // other end would not work correctly.
  always @(posedge phy_clk) begin
    if (phy_phase_valid)
      pr_phyr_tkeep_q <= {PR_phyr_tkeep[5], PR_phyr_tkeep[3], PR_phyr_tkeep[1]};
  end

  // tready will always be asserted. buffer management is handled in the RX OLLM.
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      BR_phyr_tready <= #TCQ 1'b0;
    else
      BR_phyr_tready <= #TCQ 1'b1;
  end

  // }}} ---------------------------------


  // {{{ Write Port Controller -----------
  reg [C_ADDR_LEN-1:0]  br_phy_starting_waddr;
  reg [C_ADDR_LEN-1:0]  br_phy_bram_waddr_d;

  // The write enable is simply the registered version of tready and tvalid.
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      br_phy_bram_we <= #TCQ 1'b0;
    // This is the timeout circuit! Intentionally deceptive name. Once set, it is stable, ok to be metastable.
    else if (buf_log_sof_out)
      br_phy_bram_we <= #TCQ 1'b0;
    else
      br_phy_bram_we <= #TCQ phy_phase_valid;
  end


  // Store data contiguously. Unlike the Transmit Buffer, the Receive Buffer structure
  // does not have dedicated segments for each packet. This simplifies the logic for the
  // address. However, we must briefly record the starting address for a packet in the
  // chance that the packet gets discontinued. If that happens, reload the address with
  // that stored count.
  always @* begin
    br_phy_bram_waddr_d = br_phy_bram_waddr + 1;
  end

  assign complete_packet_written = !pr_phyr_src_dsc_q && pr_phyr_tlast_q && br_phy_bram_we;
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      br_phy_starting_waddr <= #TCQ 0;
    end else if (complete_packet_written) begin
      br_phy_starting_waddr <= #TCQ br_phy_bram_waddr_d;
    end
  end
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      br_phy_bram_waddr <= #TCQ 0;
    end else if (pr_phyr_src_dsc_q && br_phy_bram_we) begin // could be qualified with pr_phyr_tlast_q
      br_phy_bram_waddr <= #TCQ br_phy_starting_waddr;
    end else if (br_phy_bram_we) begin
      br_phy_bram_waddr <= #TCQ br_phy_bram_waddr_d;
    end
  end


    // *- COVERAGE (BR_br_phy_bram_waddr_enumerate)
    // enumerate br_phy_bram_waddr crossed with RX_DEPTH

    // *- COVERAGE (BR_br_phy_bram_waddr_rollover)
    // Observe that br_phy_bram_waddr rolls over

    // *- COVERAGE (BR_br_phy_bram_waddr_cross_tlast)
    // Cross br_phy_bram_waddr with PR_phyr_tlast

    // *- COVERAGE (BR_br_phy_bram_waddr_reload)
    // Observe a discontinue event

    // *- COVERAGE (BR_complete_packet_written_b2b)
    // Observe complete_packet_written assert for two consecutive clock cycles

    // *- COVERAGE (BR_complete_packet_written_b2b2b)
    // Observe complete_packet_written assert for three consecutive clock cycles

    // *- COVERAGE (BR_reset_br_phy_starting_waddr_non_zero)
    // Observe a reset when br_phy_starting_waddr is non-zero

    // *- COVERAGE (BR_reset_br_phy_bram_waddr_non_zero)
    // Observe a reset when br_phy_bram_waddr is non-zero

  // }}} ---------------------------------


  // {{{ Write Flow Control --------------

  // keeps track of the number of free, full-sized packets the buffer is capable of storing.
  // Take the difference between the two address pointers and divide by the largest sized packet.
  // NOTE: using a 6-bit value for free_buf_packet_count is safe so long as the buffer is capable of
  // storing 64 or fewer packets. The max size for C_ADDR_LEN is 11. By shifting out 6 (C_MAX_INDEX_LEN),
  // we're left with only 5 bits. There are 6 bits because BR_phy_buf_stat is 6 bits. Since RX_DEPTH
  // can currently only be 32 max, the upper bit should be zero.
  // NOTE: free_buf_word_count won't underrun from 0 to -1 because the true size of a max packet is 34
  // though the code treats a max packet to be 64 (2^C_MAX_INDEX_LEN). So, once the buffer becomes "full"
  // there are actuall 20 (64 minus 34) free locations left.
  wire [C_ADDR_LEN-1:0] free_buf_word_count   = brp_phy_bram_raddr - br_phy_bram_waddr;
  wire [5:0]            free_buf_packet_count = (free_buf_word_count >> C_MAX_INDEX_LEN);
  wire [5:0]            br_phy_buf_stat_max;

  // Add a little bit of logic to come up with a safe value for the buf_stat.
  // special scenario for when the depth is 32:
  // A value of 31 or greater could be interpreted as rx flow control.
  // Avoid this scenario by masking anything above 30.
  // When RX_DEPTH is below 32, the logic may be simplified to not check for 30+.
  assign br_phy_buf_stat_max = (RX_DEPTH == 32) ? 6'h1E : RX_DEPTH;
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      BR_phy_buf_stat <= #TCQ br_phy_buf_stat_max;
    // raddr will sometimes roll past the waddr. This is prevents the calculation from being wrong in that case.
    end else if ((free_buf_word_count == 0) || (free_buf_word_count == 1)) begin
      BR_phy_buf_stat <= #TCQ br_phy_buf_stat_max;
    end else if (free_buf_packet_count > 30) begin
      BR_phy_buf_stat <= #TCQ br_phy_buf_stat_max;
    end else begin
      BR_phy_buf_stat <= #TCQ free_buf_packet_count;
    end
  end


    // *- COVERAGE (BR_free_buf_word_count_enumerate)
    // Enumerate free_buf_word_count

    // *- ASSERTION (BR_free_buf_word_count_range)
    // free_buf_word_count cannot fall between the range of 2 - 20

    // *- COVERAGE (BR_free_buf_packet_count_enumerate)
    // Enumerate free_buf_packet_count (0 through 32)

    // *- ASSERTION (BR_free_buf_packet_count_range)
    // free_buf_packet_count will never exceed 32

    // *- COVERAGE (BR_phy_buf_stat_enumerate)
    // Enumerate BR_phy_buf_stat (0 through 30)

    // *- ASSERTION (BR_phy_buf_stat_behavior)
    // BR_phy_buf_stat will never exceed RX_DEPTH or 30, whichever is smaller

    // *- ASSERTION (BR_phy_buf_stat_behavior)
    // BR_phy_buf_stat will never increment or decrement by more than one

    // *- COVERAGE (BR_brp_phy_bram_raddr_and_br_phy_bram_waddr_increment)
    // Observe both brp_brp_phy_bram_raddr and br_phy_bram_waddr increment on the same cycle

    // *- COVERAGE (BR_phy_buf_stat_full_then_empty)
    // Observe BR_phy_buf_stat == 30 after it once held a value of 0.

  // }}} ---------------------------------


  // {{{ BRAM Bank -----------------------
  // this will be an asynchronous FIFO when !UNIFIED_CLK.  Otherwise, it is
  // a simple synchronous FIFO/buffer.
  srio_gen2_v4_1_16_buf_rx_bram_bank
   #(.TCQ                  (TCQ),
     .UNIFIED_CLK          (UNIFIED_CLK),
     .C_FAMILY             (C_FAMILY),
     .C_ADDR_LEN           (C_ADDR_LEN))
   buf_rx_bram_bank_inst
    (.phy_clk              (phy_clk),
     .log_clk              (log_clk),
     .buf_phy_rst_q        (buf_phy_rst_q),
     .buf_log_rst_q        (buf_log_rst_q),
     // in from Physical clock
     .BR_phy_bram_waddr    (br_phy_bram_waddr),
     .BR_phy_bram_we       (br_phy_bram_we),
     .PR_phy_tdata_q       (pr_phyr_tdata_q),
     .PR_phy_tuser_q       (pr_phyr_tuser_q),
     .PR_phy_tkeep_q       (pr_phyr_tkeep_q),
     .PR_phy_tlast_q       (pr_phyr_tlast_q),
     // in/out to Logical clock
     .BR_log_bram_raddr    (br_log_bram_raddr),
     .BR_log_bram_rd       (br_log_bram_rd),
     .BRB_log_bram_tdata   (brb_log_bram_tdata),
     .BRB_log_bram_tuser   (brb_log_bram_tuser),
     .BRB_log_bram_tkeep   (brb_log_bram_tkeep),
     .BRB_log_bram_tlast   (brb_log_bram_tlast)
    );
  // }}} ---------------------------------


  // {{{ Async Passage -------------------

  // On the ports, it takes in binary values and outputs binary values.
  // Internally, this module passes Gray Coded count values between the clock domains.
  generate if (!UNIFIED_CLK) begin: async_passage_gen
    srio_gen2_v4_1_16_buf_rx_async_passage
     #(.TCQ                     (TCQ),
       .C_ADDR_LEN              (C_ADDR_LEN))
     buf_rx_async_passage_inst
      (.log_clk                 (log_clk),
       .phy_clk                 (phy_clk),
       .buf_log_rst_q           (buf_log_rst_q),
       .buf_phy_rst_q           (buf_phy_rst_q),
       .BR_log_bram_raddr       (br_log_bram_raddr),
       .BR_phy_starting_waddr   (br_phy_starting_waddr),
       .BRP_phy_bram_raddr      (brp_phy_bram_raddr),
       .BRP_log_starting_waddr  (brp_log_starting_waddr)
    );

  // when a common clock structure is used, save resources by just passing the values across
  end else                   begin: sync_passage_gen
    assign brp_phy_bram_raddr      = br_log_bram_raddr;
    assign brp_log_starting_waddr  = br_phy_starting_waddr;

  end
  endgenerate


    // *- COVERAGE (BR_brp_phy_bram_raddr_jumps_by_2)
    // Observe that brp_phy_bram_raddr increments by 2

    // *- COVERAGE (BR_brp_phy_bram_raddr_jumps_by_3)
    // Observe that brp_phy_bram_raddr increments by 3

    // *- COVERAGE (BR_brp_phy_bram_raddr_jumps_by_4)
    // Observe that brp_phy_bram_raddr increments by 4

    // *- COVERAGE (BR_brp_log_starting_waddr_jumps_by_2)
    // Observe that brp_log_starting_waddr increments by 2

    // *- COVERAGE (BR_brp_log_starting_waddr_jumps_by_3)
    // Observe that brp_log_starting_waddr increments by 3

    // *- COVERAGE (BR_brp_log_starting_waddr_jumps_by_4)
    // Observe that brp_log_starting_waddr increments by 4

  // }}} ---------------------------------

 
  // {{{ Read Flow Control ---------------

  wire [C_ADDR_LEN-1:0]  log_count_diff = brp_log_starting_waddr - br_log_bram_raddr;
  wire                   last_present_d = brb_log_bram_tlast && 
                                          // conditions by which we advance the final pipeline stage -
                                          ((BR_bufr_tvalid && LE_bufr_tready) ||
                                          (br_bufr_tvalid_d[1] && !BR_bufr_tvalid));


  // The buffer empty signal should assert at the end of the packet that makes it go empty.
  // If the buffer goes empty, the logic was designed to specifically make sure the empty signal
  // doesn't clear until the previous packet has completely pushed through the pipeline. This
  // can be observed by the addition of tvalid and tvalid_q on log_clr_empty
  assign log_set_empty  = log_set_empty_condition && last_present_d && !log_buffer_empty;
  assign log_clr_empty  = (log_count_diff != 0) && !br_bufr_tvalid_q && !BR_bufr_tvalid;
  always @(posedge log_clk) begin
    if (buf_log_rst_q)
      log_buffer_empty <= #TCQ 1'b1;
    else if (log_set_empty)
      log_buffer_empty <= #TCQ 1'b1;
    else if (log_clr_empty)
      log_buffer_empty <= #TCQ 1'b0;
  end

  always @(posedge log_clk) begin
    if (log_count_diff == 0)
      log_set_empty_condition <= #TCQ 1'b1;
    else if (log_clr_empty)
      log_set_empty_condition <= #TCQ 1'b0;
  end


    // *- COVERAGE (BR_log_set_empty_and_log_clr_empty)
    // log_set_empty and log_clr_empty are expected to occasionally overlap. Observe this event.

  // }}} ---------------------------------


  // {{{ Read Port Controller ------------

  assign br_log_bram_rd       = (log_pipeline_vacancy || (BR_bufr_tvalid && LE_bufr_tready)) && !log_buffer_empty;
  assign log_pipeline_vacancy = log_pipeline_count < 3 ? 1 : 0;

  // There are 3 stages of pipeline between the buffer and the interface. As a result,
  // we must keep track of a counter that tells how many data beats are sitting between
  // the buffer and the interface. i.e. how many stages of the pipeline are full.
  always @(posedge log_clk) begin
    if (buf_log_rst_q)
      log_pipeline_count <= #TCQ 2'h0;
    else if (log_buffer_empty)
      log_pipeline_count <= #TCQ 2'h0;
    else if (br_log_bram_rd && !(BR_bufr_tvalid && LE_bufr_tready))
      log_pipeline_count <= #TCQ log_pipeline_count + 1;
  end

  // This is a contiguous address. There are no gaps between packets in the memory. As a
  // result, simply increment when data is captured. When the buffer becomes empty, subtract
  // by one. This is done in order to close up the final packet on empty and prepare for
  // the next packet when the buffer becomes unempty.
  // Add a bit of abstraction here with the _op signal in order to make sure the tools don't
  // infer two adders when only one is needed.
  wire [C_ADDR_LEN-1:0] br_log_bram_raddr_op = log_set_empty ? -1 : 1;
  always @(posedge log_clk) begin
    if (buf_log_rst_q) begin
      br_log_bram_raddr <= #TCQ 0;
    end else if (log_set_empty) begin
      br_log_bram_raddr <= #TCQ br_log_bram_raddr + br_log_bram_raddr_op;
    end else if (br_log_bram_rd) begin
      br_log_bram_raddr <= #TCQ br_log_bram_raddr + br_log_bram_raddr_op;
    end
  end


    // *- COVERAGE (BR_br_log_bram_raddr_enumerate)
    // Enumerate br_log_bram_raddr crossed with RX_DEPTH

    // *- COVERAGE (BR_br_log_bram_raddr_rollover)
    // Observe br_log_bram_raddr rolls over

    // *- ASSERTION (BR_log_pipeline_count_behavior)
    // log_pipeline_count never wraps (3 -> 0) except on log_buffer_empty

    // *- COVERAGE (BR_br_log_bram_raddr_cross_tlast)
    // Cross br_log_bram_raddr with BR_bufr_tlast

    // *- COVERAGE (BR_reset_br_log_bram_raddr_non_zero)
    // Observe a reset when br_log_bram_raddr is non-zero

    // *- COVERAGE (BR_log_pipeline_count_transitions)
    // Observe the following transitions on log_pipeline_count:
    // 0 -> 1, 1 -> 2, 2 -> 3, 3 -> 2, 2-> 1, 1 -> 0
    // and when the buffer goes empty: 3 -> 0, 2 -> 0

  // }}} ---------------------------------


  // {{{ LOG Interface -------------------

  // advance the pipeline if the log layer is ready or if the
  // buffer does not currently have anything valid on the bus
  reg buf_tstart_q;
  wire bufr_advance_condition = LE_bufr_tready || !BR_bufr_tvalid;


  // TLAST generation -
  // hold tlast if the logical layer's tready is not asserted. Otherwise,
  // take the next value.
  always @(posedge log_clk) begin
    if (buf_log_rst_q) begin
      BR_bufr_tlast <= #TCQ 1'b0;
    end else if (bufr_advance_condition) begin
      // NOTE: advancing the control signals can be tricky
      // for simplification, here are the conditions under which we enter this case:
      // TREADY = 0, TVALID = 0, tvalid_d = 1
      // TREADY = 1, TVALID = 0, tvalid_d = 1
      // TREADY = 1, TVALID = 1, tvalid_d = x
      if (br_bufr_tvalid_d[1] || BR_bufr_tvalid)
        BR_bufr_tlast <= #TCQ brb_log_bram_tlast;
    end
  end

  // TSTART generation -
  // This is not part of the AXI specification but is a very useful signal
  // It gets passed through the TUSER bus.
  // NOTE: This signal was specifically created to ease timing in the LOG
  always @* begin
    buf_tstart = buf_tstart_q;
    if (BR_bufr_tlast && (LE_bufr_tready && BR_bufr_tvalid)) begin
      buf_tstart = 1'b1;
    end else if (LE_bufr_tready && BR_bufr_tvalid) begin
      buf_tstart = 1'b0;
    end
  end
  always @(posedge log_clk) begin
    if (buf_log_rst_q) begin
      buf_tstart_q <= #TCQ 1'b1;
    end else begin
      buf_tstart_q <= #TCQ buf_tstart;
    end
  end

  // general bufr signal generation
  // register outgoing data fields. Since this is going to the user, add a reset.
  always @(posedge log_clk) begin
    if (buf_log_rst_q) begin
      BR_bufr_tdata  <= #TCQ 64'h0;
      BR_bufr_tuser  <= #TCQ 8'h0;
      BR_bufr_tvalid <= #TCQ 1'b0;
    end else if (bufr_advance_condition) begin
      BR_bufr_tdata  <= #TCQ brb_log_bram_tdata;
      BR_bufr_tuser  <= #TCQ {4'h0, buf_tstart, brb_log_bram_tuser, 1'b0};
      BR_bufr_tvalid <= #TCQ (br_bufr_tvalid_d[1] || BR_bufr_tvalid) && !log_buffer_empty;
    end
  end


  // TSTRB generation/reconstruction -
  // convert the simplified internal strobe value back to its 8-bit value.
  // If more combinations of strobe become acceptable, this will take a redesign.
  always @(posedge log_clk) begin
    if (buf_log_rst_q) begin
      BR_bufr_tkeep <= #TCQ 8'h0;
    end else if (bufr_advance_condition) begin
      if (!brb_log_bram_tlast)
        BR_bufr_tkeep <= #TCQ 8'hFF;
      else
        BR_bufr_tkeep <= #TCQ {1'b0, brb_log_bram_tkeep[2], brb_log_bram_tkeep[2], brb_log_bram_tkeep[1], 
                               brb_log_bram_tkeep[1], brb_log_bram_tkeep[0], brb_log_bram_tkeep[0], 1'b1};
    end
  end


  // pipeline TVALID generation -
  always @(posedge log_clk) begin
    if (buf_log_rst_q) begin
      br_bufr_tvalid_d <= #TCQ 2'b0;
      br_bufr_tvalid_q <= #TCQ 1'b0;
    end else begin
      br_bufr_tvalid_d <= #TCQ {br_bufr_tvalid_d[0], br_log_bram_rd};
      br_bufr_tvalid_q     <= #TCQ BR_bufr_tvalid;
    end
  end

  // }}} ---------------------------------


  // {{{ EVAL timer ----------------------
  // the signal names in the following code are deliberately vague and
  // misleading.  When the eval parameter is selected, this unit will be
  // present.  When the timer expires, buf_log_sof_out will assert to 1, and not
  // release until a reset.
  generate if (EVAL) begin: lnk_sof_gen
    reg [7:0] log_sof_clr = 8'hFF;
    always @(posedge log_clk) begin
      log_sof_clr <= #TCQ {log_sof_clr[6:0], 1'b0};
    end

    // FIXME - CFR - take into account MODE_XG
    srio_gen2_v4_1_16_eval sof_gen_inst
     (.ena      (1'b1),
      .x        (buf_log_sof_out_d),
      .pci_rst  (log_sof_clr[7]),
      .pci_clk  (log_clk)
     );

  end else           begin: lnk_sof_gen

    assign buf_log_sof_out_d = 1'b0;

  end
  endgenerate
  always @(posedge log_clk) begin
    buf_log_sof_out <= #TCQ buf_log_sof_out_d;
  end

  // }}} ---------------------------------


endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/buf/srio_gen2_v4_1_16_buf_rx_async_passage.v#1 $
//
// BUF_RX_ASYNC_PASSAGE
// Description:
// This module allows the passage of information between the physical
// and logical clock domains.
//   
// Hierarchy:
// BUF_TOP
//  |______BUF_TX
//  |____________BUF_TX_SYNC_UNIT
//  |____________BUF_TX_BRAM_BANK
//  |______BUF_RX
//  |____________BUF_RX_ASYNC_PASSAGE <-- this module
//  |____________BUF_RX_BRAM_BANK
//----------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)

module srio_gen2_v4_1_16_buf_rx_async_passage
  #(
    parameter TCQ           = 100,
    parameter C_ADDR_LEN    = 11)                        // {11, 12, 13}
   (
   // {{{ port declarations ----------------- 
    input                       log_clk,                 // Freerunning Logical Layer clk
    input                       phy_clk,                 // Freerunning Physical Layer clk
    input                       buf_log_rst_q,           // Synchronous Logical Layer rst
    input                       buf_phy_rst_q,           // Synchronous Physical Layer rst
    // Signals to/from the RX Buffer
    input      [C_ADDR_LEN-1:0] BR_log_bram_raddr,       // read address from log domain
    input      [C_ADDR_LEN-1:0] BR_phy_starting_waddr,   // write packet count from phy domain
    output reg [C_ADDR_LEN-1:0] BRP_phy_bram_raddr,      // read address ported to phy domain
    output reg [C_ADDR_LEN-1:0] BRP_log_starting_waddr   // write packet count ported to log domain
   // }}} --------------------------------- 
   );


  // {{{ wire declarations ---------------

  // signals for converting the read address
  reg  [C_ADDR_LEN-1:0]  log_bram_raddr_gc;           // Gray code for the read address
  (* ASYNC_REG = "TRUE" *)
  reg  [C_ADDR_LEN-1:0]  phy_bram_raddr_gc_async;     // first capture of read address in phy domain
  reg  [C_ADDR_LEN-1:0]  phy_bram_raddr_gc;           // second capture of read address in phy domain
  reg  [C_ADDR_LEN-1:0]  brp_phy_bram_raddr_d;        // combinatorial transform of Gray to binary of read address

  // signals for converting the starting write address
  reg  [C_ADDR_LEN-1:0]  phy_starting_waddr_gc;       // Gray code for the write packet
  (* ASYNC_REG = "TRUE" *)
  reg  [C_ADDR_LEN-1:0]  log_starting_waddr_gc_async; // first capture of write packet in log domain
  reg  [C_ADDR_LEN-1:0]  log_starting_waddr_gc;       // second capture of write packet in log domain
  reg  [C_ADDR_LEN-1:0]  brp_log_starting_waddr_d;    // combinatorial transform of Gray to binary of write packet

  // }}} ---------------------------------


  // {{{ Functions -----------------------

  // Gray Code works by XORing consecutive bits together. For a 4-bit conversion:
  // GrayCode[0] = BinaryCode[0] ^ BinaryCode[1]
  // GrayCode[1] = BinaryCode[1] ^ BinaryCode[2]
  // GrayCode[2] = BinaryCode[2] ^ BinaryCode[3]
  // GrayCode[3] = BinaryCode[3]
  function [C_ADDR_LEN-1:0] binary_to_gray_code(input [C_ADDR_LEN-1:0] binary_value);
  begin
      binary_to_gray_code = (binary_value >> 1) ^ binary_value;
  end
  endfunction

  // Conversion back to Binary is the reverse of the procedure to convert to Gray. For a 4-bit conversion:
  // BinaryCode[3] = GrayCode[3]
  // BinaryCode[2] = GrayCode[2] ^ BinaryCode[3]
  // BinaryCode[1] = GrayCode[1] ^ BinaryCode[2]
  // BinaryCode[0] = GrayCode[0] ^ BinaryCode[1]
  function [C_ADDR_LEN-1:0] gray_code_to_binary(input [C_ADDR_LEN-1:0] gray_value);
  begin : gray_code_to_binary_logic
      integer xx;

      for (xx = 0; xx < C_ADDR_LEN; xx = xx + 1) begin
          gray_code_to_binary[xx] = ^(gray_value >> xx);
      end
  end
  endfunction

  // }}} ---------------------------------


  // BRP_phy_bram_raddr generation -
  // Use Gray coding when the clocks aren't synchronized to pass tags between
  // the two domains.

  // {{{ BR_log_bram_raddr passing -------

  // convert the binary value of the read address to Gray
  always @(posedge log_clk) begin
    if (buf_log_rst_q)
      log_bram_raddr_gc <= #TCQ 0;
    else
      log_bram_raddr_gc <= #TCQ binary_to_gray_code(BR_log_bram_raddr);
  end


  // synchronizing registers. Since only one bit changes per transition, 
  // simply double-registering is sufficient.
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q) begin
      phy_bram_raddr_gc_async <= #TCQ 0;
      phy_bram_raddr_gc       <= #TCQ 0;
    end else begin
      phy_bram_raddr_gc_async <= #TCQ log_bram_raddr_gc;
      phy_bram_raddr_gc       <= #TCQ phy_bram_raddr_gc_async;
    end
  end


  // convert the read address Gray Code back to binary
  always @* begin
    brp_phy_bram_raddr_d = gray_code_to_binary(phy_bram_raddr_gc);
  end


  // Final register of the read address.
  // For those of you keeping track, it takes 1 log_clk cycle and 3 phy_clk cycles to transfer the address
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      BRP_phy_bram_raddr <= #TCQ 0;
    else
      BRP_phy_bram_raddr <= #TCQ brp_phy_bram_raddr_d;
  end


    // *- COVERAGE (BR_phy_bram_raddr_gc_enumerate)
    // Enumerate phy_bram_raddr_gc

  // }}} ---------------------------------

  // End BRP_phy_bram_raddr generation


  // BRP_log_starting_waddr generation -
  // Use Gray coding when the clocks aren't synchronized to pass tags between
  // the two domains.

  // {{{ BR_phy_starting_waddr passing -------

  // convert the binary value of the starting write address to Gray
  always @(posedge phy_clk) begin
    if (buf_phy_rst_q)
      phy_starting_waddr_gc <= #TCQ 0;
    else
      phy_starting_waddr_gc <= #TCQ binary_to_gray_code(BR_phy_starting_waddr);
  end


  // synchronizing registers. Since only one bit changes per transition, 
  // simply double-registering is sufficient.
  always @(posedge log_clk) begin
    if (buf_log_rst_q) begin
      log_starting_waddr_gc_async <= #TCQ 0;
      log_starting_waddr_gc       <= #TCQ 0;
    end else begin
      log_starting_waddr_gc_async <= #TCQ phy_starting_waddr_gc;
      log_starting_waddr_gc       <= #TCQ log_starting_waddr_gc_async;
    end
  end


  // convert the read address Gray Code back to binary
  always @* begin
    brp_log_starting_waddr_d = gray_code_to_binary(log_starting_waddr_gc);
  end


  // Final register of the starting write address.
  // For those of you keeping track, it takes 1 phy_clk cycle and 3 log_clk cycles to transfer the address
  always @(posedge log_clk) begin
    if (buf_log_rst_q)
      BRP_log_starting_waddr <= #TCQ 0;
    else
      BRP_log_starting_waddr <= #TCQ brp_log_starting_waddr_d;
  end


    // *- COVERAGE (BR_phy_starting_waddr_gc_enumerate)
    // Enumerate phy_starting_waddr_gc

  // }}} ---------------------------------

  // End BRP_log_starting_waddr generation

endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/buf/srio_gen2_v4_1_16_eval.v#1 $
//----------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)

module srio_gen2_v4_1_16_eval
#(parameter TCQ = 100)
(
                ena,
                x,
                pci_rst,
                pci_clk
                );


  // Declare the port directions.

  input         ena;
  output        x;
  input         pci_rst;
  input         pci_clk;


  //******************************************************************//
  // Stage A.                                                         //
  //******************************************************************//


  reg     [7:0] a = 8'h00;
  reg           a_out = 1'b0;
  wire          a_ceo;
  wire          a_en;

  assign a_en = 1'b1;

  always @(posedge pci_clk or posedge pci_rst) begin : xpci_a
    if (pci_rst) begin
      a <= #TCQ 8'h00;
      a_out <= #TCQ 1'b0;
    end else begin
      if (a_en) begin
        a <= #TCQ a + 8'h01;
      end
      a_out <= #TCQ a_ceo;
    end
  end

  assign a_ceo = a_en & (a == 8'hff);


  //******************************************************************//
  // Stage B.                                                         //
  //******************************************************************//


  reg     [7:0] b = 8'h00;
  reg           b_out = 1'b0;
  wire          b_ceo;
  wire          b_en;

  assign b_en = a_out;

  always @(posedge pci_clk or posedge pci_rst) begin : xpci_b
    if (pci_rst) begin
      b <= #TCQ 8'h00;
      b_out <= #TCQ 1'b0;
    end else begin
      if (b_en) begin
        b <= #TCQ b + 8'h01;
      end
      b_out <= #TCQ b_ceo;
    end
  end

  assign b_ceo = b_en & (b == 8'hff);


  //******************************************************************//
  // Stage C.                                                         //
  //******************************************************************//


  reg     [7:0] c = 8'h00;
  reg           c_out = 1'b0;
  wire          c_ceo;
  wire          c_en;

  assign c_en = b_out;

  always @(posedge pci_clk or posedge pci_rst) begin : xpci_c
    if (pci_rst) begin
      c <= #TCQ 8'h00;
      c_out <= #TCQ 1'b0;
    end else begin
      if (c_en) begin
        c <= #TCQ c + 8'h01;
      end
      c_out <= #TCQ c_ceo;
    end
  end

  assign c_ceo = c_en & (c == 8'hff);


  //******************************************************************//
  // Stage D.                                                         //
  //******************************************************************//


  reg     [7:0] d = 8'h00;
  reg           d_out = 1'b0;
  wire          d_ceo;
  wire          d_en;

  assign d_en = c_out;

  always @(posedge pci_clk or posedge pci_rst) begin : xpci_d
    if (pci_rst) begin
      d <= #TCQ 8'h00;
      d_out <= #TCQ 1'b0;
    end else begin
      if (d_en) begin
        d <= #TCQ d + 8'h01;
      end
      d_out <= #TCQ d_ceo;
    end
  end

  assign d_ceo = d_en & (d == 8'hff);


  //******************************************************************//
  // Stage E.                                                         //
  //******************************************************************//


  reg     [7:0] e = 8'h00;
  wire          e_ceo;
  wire          e_en;

  assign e_en = d_out;

  always @(posedge pci_clk or posedge pci_rst) begin : xpci_e
    if (pci_rst) begin
      e <= #TCQ 8'h00;
    end else begin
      if (e_en) begin
        e <= #TCQ e + 8'h01;
      end
    end
  end

  assign e_ceo = e_en & (e == 8'hff);


  //******************************************************************//
  // Generate the expire flag.                                        //
  //******************************************************************//


  reg           bug_fix = 1'b0;

  always @(posedge pci_clk or posedge pci_rst) begin : xpci_bug_fix
    if (pci_rst)
      bug_fix <= #TCQ 1'b0;
    else if (e_ceo)
      bug_fix <= #TCQ 1'b1;
  end

  assign x = bug_fix & ena;


  //******************************************************************//
  //                                                                  //
  //******************************************************************//


endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/buf/srio_gen2_v4_1_16_buf_tx_sync_unit.v#4 $
//----------------------------------------------------------------------
//
// BUF_TX_SYNC_UNIT
// Description:
// This module facilitates the passage of packet data from the logical
// clock domain to the physical clock domain.
//
// Hierarchy:
// BUF_TOP
//  |______BUF_TX
//  |____________BUF_TX_SYNC_UNIT <-- this module
//  |____________BUF_TX_BRAM_BANK
//  |______BUF_RX
//  |____________BUF_RX_ASYNC_PASSAGE
//  |____________BUF_RX_BRAM_BANK
`timescale 1ps/1ps

module srio_gen2_v4_1_16_buf_tx_sync_unit
  #(
    parameter TCQ           = 100,
    parameter C_FAMILY      = "virtex6",     // {virtex5, virtex6, virtex7, spartan6, spartan7}
    parameter TX_DEPTH      = 8,             // {8, 16, 32}
    parameter UNIFIED_CLK   = 0)             // {0, 1}
   (
   // {{{ port declarations -----------------

    input             log_clk,               // Freerunning Logical Layer clock
    input             phy_clk,               // Freerunning Physical Layer clock
    input             buf_log_rst_q,         // Synchronous Logical Layer reset
    input             buf_phy_rst_q,         // Synchronous Physical Layer reset
    // LOG TX Interface
    input             LD_buft_tlast,         // Last Beat
    input             LD_buft_tvalid,        // Valid Packet Beat
    output reg        BTS_buft_tready,       // Packet Beat Accepted
    input   [7:0]     LD_buft_tkeep,         // Valid Bytes in this beat, only valid on last
    input   [63:0]    LD_buft_tdata,         // Packet Data
    input   [7:0]     LD_buft_tuser,         // {3'h0, Response, 1'b0, VC, CRF, 1'b0} AXI Compliance Pad
    output reg        BTS_response_only,     // Buffer only has room for Resp Packets
    // PHY clock domain signals
    input             PC_master_enable,      // Master Enable Indication
    output [63:0]     BTS_tx_data,           // Data Out
    output            BTS_tx_start,          // Start of Frame
    output            BTS_tx_last,           // End of Frame
    output            BTS_tx_valid,          // Source Data Ready
    output [7:0]      BTS_tx_user,           // Critical Request Flow
    output [2:0]      BTS_tx_keep,           // Remainder
    input             BT_tx_ready,           // Destination Data Ready
    input             BT_packet_ack          // Packet Accepted Intication

   // }}} ---------------------------------
   );

  // {{{ local parameters ------------------

    // dial this value in for more or less buffer space dedicated to responses
  localparam RESPONSE_ONLY_THRESHOLD = 2;
  localparam PTR_WIDTH = TX_DEPTH == 8  ? 3 :
                         TX_DEPTH == 16 ? 4 : 5;
  // }}} ---------------------------------


  // {{{ wire declarations -----------------
  reg  [5:0] outstanding_packets;     // there is at least 1 more bit than TX_DEPTH because we can capture more packets
  wire       log_packet_available_n;  // indicates when a packet has been released
  wire       outstanding_packets_inc; // + 1 to outstanding packets
  wire       outstanding_packets_dec; // - 1 to outstanding packets
  reg        pcfg_master_en_a;        // synchronization registers
  reg        bts_buft_tstart;         // sop signal made to look like an AXI signal
  wire       afifo_full;              // full indication - only req'd for real_sync_unit but used in coverage


    // *- COVERAGE (BT_outstanding_packets_enumerate)
    // Enumerate outstanding_packets across all valid values (0 through TX_DEPTH + 16)

    // *- ASSERTION (BT_outstanding_packets_behavior)
    // outstanding packets never increments or decrements by more that 1.

    // *- COVERAGE (BT_outstanding_packets_inc_dec)
    // Show that both the increment and decrement condition happen on the same cycle

    // *- COVERAGE (BT_observe_afifo_full)
    // See that the synchronization buffer goes full.

  // }}} -----------------------------------

  generate if (!UNIFIED_CLK) begin: real_sync_unit
    // {{{ Real Synch Unit ---

    // we only use these signals when the dist ram is instantiated - no need to
    // create them otherwise.
    wire        afifo_empty;
    wire [71:0] afifo_rdata;
    wire        afifo_rd    = BT_tx_ready;
    wire        afifo_wr    = LD_buft_tvalid && BTS_buft_tready;
    wire [71:0] afifo_wdata = {bts_buft_tstart, LD_buft_tlast,
                               LD_buft_tkeep[5], LD_buft_tkeep[3], LD_buft_tkeep[1],
                               LD_buft_tuser[2:1], LD_buft_tuser[4], LD_buft_tdata};


      assign BTS_tx_valid     = !afifo_empty;
      assign BTS_tx_start     = afifo_rdata[71];
      assign BTS_tx_last      = afifo_rdata[70];
      assign BTS_tx_keep      = afifo_rdata[69:67];
      assign BTS_tx_user      = {3'h0, afifo_rdata[64], 1'b0, afifo_rdata[66:65], 1'b0};
      assign BTS_tx_data      = afifo_rdata[63:0];

      always @(posedge log_clk) begin
        if (buf_log_rst_q)
          BTS_buft_tready <= #TCQ 1'b0;
        else
          BTS_buft_tready <= !afifo_full;
      end

    fifo_generator_vlog_beh
     // {{{ parameter list ---------------
     #(.C_COMMON_CLOCK                 (0),
       .C_COUNT_TYPE                   (0),
       .C_DATA_COUNT_WIDTH             (4),
       .C_DEFAULT_VALUE                ("BlankString"),
       .C_DIN_WIDTH                    (72),
       .C_DOUT_RST_VAL                 ("0"),
       .C_DOUT_WIDTH                   (72),
       .C_ENABLE_RLOCS                 (0),
       .C_ENABLE_RST_SYNC              (1),
       .C_ERROR_INJECTION_TYPE         (0),
       .C_FAMILY                       (C_FAMILY),
       .C_FULL_FLAGS_RST_VAL           (1),
       .C_HAS_ALMOST_EMPTY             (0),
       .C_HAS_ALMOST_FULL              (1),
       .C_HAS_BACKUP                   (0),
       .C_HAS_DATA_COUNT               (0),
       .C_HAS_INT_CLK                  (0),
       .C_HAS_MEMINIT_FILE             (0),
       .C_HAS_OVERFLOW                 (0),
       .C_HAS_RD_DATA_COUNT            (0),
       .C_HAS_RD_RST                   (0),
       .C_HAS_RST                      (1),
       .C_HAS_SRST                     (0),
       .C_HAS_UNDERFLOW                (0),
       .C_HAS_VALID                    (0),
       .C_HAS_WR_ACK                   (0),
       .C_HAS_WR_DATA_COUNT            (0),
       .C_HAS_WR_RST                   (0),
       .C_IMPLEMENTATION_TYPE          (2),
       .C_INIT_WR_PNTR_VAL             (0),
       .C_MEMORY_TYPE                  (2),
       .C_MIF_FILE_NAME                ("BlankString"),
       .C_MSGON_VAL                    (1),
       .C_OPTIMIZATION_MODE            (0),
       .C_OVERFLOW_LOW                 (0),
       .C_PRELOAD_LATENCY              (0),
       .C_PRELOAD_REGS                 (1),
       .C_PRIM_FIFO_TYPE               ("512x72"),
       .C_PROG_EMPTY_THRESH_ASSERT_VAL (4),
       .C_PROG_EMPTY_THRESH_NEGATE_VAL (5),
       .C_PROG_EMPTY_TYPE              (0),
       .C_PROG_FULL_THRESH_ASSERT_VAL  (13),
       .C_PROG_FULL_THRESH_NEGATE_VAL  (12),
       .C_PROG_FULL_TYPE               (0),
       .C_RD_DATA_COUNT_WIDTH          (4),
       .C_RD_DEPTH                     (16),
       .C_RD_FREQ                      (1),
       .C_RD_PNTR_WIDTH                (4),
       .C_UNDERFLOW_LOW                (0),
       .C_USE_DOUT_RST                 (1),
       .C_USE_ECC                      (0),
       .C_USE_EMBEDDED_REG             (0),
       .C_USE_FIFO16_FLAGS             (0),
       .C_USE_FWFT_DATA_COUNT          (0),
       .C_VALID_LOW                    (0),
       .C_WR_ACK_LOW                   (0),
       .C_WR_DATA_COUNT_WIDTH          (4),
       .C_WR_DEPTH                     (16),
       .C_WR_FREQ                      (1),
       .C_WR_PNTR_WIDTH                (4),
       .C_WR_RESPONSE_LATENCY          (1),
       
       //--- below parameters are newly added in v12_0, left default
       .C_POWER_SAVING_MODE		(0),        
       .C_SYNCHRONIZER_STAGE		(2),        
       .C_INTERFACE_TYPE		(0),        
       .C_AXI_TYPE			(1),        
       .C_HAS_AXI_WR_CHANNEL		(1),        
       .C_HAS_AXI_RD_CHANNEL		(1),        
       .C_HAS_SLAVE_CE			(0),        
       .C_HAS_MASTER_CE			(0),        
       .C_ADD_NGC_CONSTRAINT		(0),        
       .C_USE_COMMON_OVERFLOW		(0),        
       .C_USE_COMMON_UNDERFLOW		(0),        
       .C_USE_DEFAULT_SETTINGS		(0),        
       .C_AXI_ID_WIDTH			(1),        
       .C_AXI_ADDR_WIDTH		(32),       
       .C_AXI_DATA_WIDTH		(64),       
       .C_AXI_LEN_WIDTH			(8),        
       .C_AXI_LOCK_WIDTH		(1),        
       .C_HAS_AXI_ID			(0),        
       .C_HAS_AXI_AWUSER		(0),        
       .C_HAS_AXI_WUSER			(0),        
       .C_HAS_AXI_BUSER			(0),        
       .C_HAS_AXI_ARUSER		(0),        
       .C_HAS_AXI_RUSER			(0),        
       .C_AXI_ARUSER_WIDTH		(1),        
       .C_AXI_AWUSER_WIDTH		(1),        
       .C_AXI_WUSER_WIDTH		(1),        
       .C_AXI_BUSER_WIDTH		(1),        
       .C_AXI_RUSER_WIDTH		(1),        
       .C_HAS_AXIS_TDATA		(1),        
       .C_HAS_AXIS_TID			(0),        
       .C_HAS_AXIS_TDEST		(0),        
       .C_HAS_AXIS_TUSER		(1),        
       .C_HAS_AXIS_TREADY		(1),        
       .C_HAS_AXIS_TLAST		(0),        
       .C_HAS_AXIS_TSTRB		(0),        
       .C_HAS_AXIS_TKEEP		(0),        
       .C_AXIS_TDATA_WIDTH		(8),        
       .C_AXIS_TID_WIDTH		(1),        
       .C_AXIS_TDEST_WIDTH		(1),        
       .C_AXIS_TUSER_WIDTH		(4),        
       .C_AXIS_TSTRB_WIDTH		(1),        
       .C_AXIS_TKEEP_WIDTH		(1),        
       .C_WACH_TYPE			(0),        
       .C_WDCH_TYPE			(0),        
       .C_WRCH_TYPE			(0),        
       .C_RACH_TYPE			(0),        
       .C_RDCH_TYPE			(0),        
       .C_AXIS_TYPE			(0),        
       .C_IMPLEMENTATION_TYPE_WACH	(1),        
       .C_IMPLEMENTATION_TYPE_WDCH	(1),        
       .C_IMPLEMENTATION_TYPE_WRCH	(1),        
       .C_IMPLEMENTATION_TYPE_RACH	(1),        
       .C_IMPLEMENTATION_TYPE_RDCH	(1),        
       .C_IMPLEMENTATION_TYPE_AXIS	(1),        
       .C_APPLICATION_TYPE_WACH		(0),        
       .C_APPLICATION_TYPE_WDCH		(0),        
       .C_APPLICATION_TYPE_WRCH		(0),        
       .C_APPLICATION_TYPE_RACH		(0),        
       .C_APPLICATION_TYPE_RDCH		(0),        
       .C_APPLICATION_TYPE_AXIS		(0),        
       .C_PRIM_FIFO_TYPE_WACH		("512x36"), 
       .C_PRIM_FIFO_TYPE_WDCH		("1kx36"),  
       .C_PRIM_FIFO_TYPE_WRCH		("512x36"), 
       .C_PRIM_FIFO_TYPE_RACH		("512x36"), 
       .C_PRIM_FIFO_TYPE_RDCH		("1kx36"),  
       .C_PRIM_FIFO_TYPE_AXIS		("1kx18"),  
       .C_USE_ECC_WACH			(0),        
       .C_USE_ECC_WDCH			(0),        
       .C_USE_ECC_WRCH			(0),        
       .C_USE_ECC_RACH			(0),        
       .C_USE_ECC_RDCH			(0),        
       .C_USE_ECC_AXIS			(0),        
       .C_ERROR_INJECTION_TYPE_WACH	(0),        
       .C_ERROR_INJECTION_TYPE_WDCH	(0),        
       .C_ERROR_INJECTION_TYPE_WRCH	(0),        
       .C_ERROR_INJECTION_TYPE_RACH	(0),        
       .C_ERROR_INJECTION_TYPE_RDCH	(0),        
       .C_ERROR_INJECTION_TYPE_AXIS	(0),        
       .C_DIN_WIDTH_WACH		(32),       
       .C_DIN_WIDTH_WDCH		(64),       
       .C_DIN_WIDTH_WRCH		(2),        
       .C_DIN_WIDTH_RACH		(32),       
       .C_DIN_WIDTH_RDCH		(64),       
       .C_DIN_WIDTH_AXIS		(1),        
       .C_WR_DEPTH_WACH			(16),       
       .C_WR_DEPTH_WDCH			(1024),     
       .C_WR_DEPTH_WRCH			(16),       
       .C_WR_DEPTH_RACH			(16),       
       .C_WR_DEPTH_RDCH			(1024),     
       .C_WR_DEPTH_AXIS			(1024),     
       .C_WR_PNTR_WIDTH_WACH		(4),        
       .C_WR_PNTR_WIDTH_WDCH		(10),       
       .C_WR_PNTR_WIDTH_WRCH		(4),        
       .C_WR_PNTR_WIDTH_RACH		(4),        
       .C_WR_PNTR_WIDTH_RDCH		(10),       
       .C_WR_PNTR_WIDTH_AXIS		(10),       
       .C_HAS_DATA_COUNTS_WACH		(0),        
       .C_HAS_DATA_COUNTS_WDCH		(0),        
       .C_HAS_DATA_COUNTS_WRCH		(0),        
       .C_HAS_DATA_COUNTS_RACH		(0),        
       .C_HAS_DATA_COUNTS_RDCH		(0),        
       .C_HAS_DATA_COUNTS_AXIS		(0),        
       .C_HAS_PROG_FLAGS_WACH		(0),        
       .C_HAS_PROG_FLAGS_WDCH		(0),        
       .C_HAS_PROG_FLAGS_WRCH		(0),        
       .C_HAS_PROG_FLAGS_RACH		(0),        
       .C_HAS_PROG_FLAGS_RDCH		(0),        
       .C_HAS_PROG_FLAGS_AXIS		(0),        
       .C_PROG_FULL_TYPE_WACH		(0),        
       .C_PROG_FULL_TYPE_WDCH		(0),        
       .C_PROG_FULL_TYPE_WRCH		(0),        
       .C_PROG_FULL_TYPE_RACH		(0),        
       .C_PROG_FULL_TYPE_RDCH		(0),        
       .C_PROG_FULL_TYPE_AXIS		(0),        
       .C_PROG_FULL_THRESH_ASSERT_VAL_WACH (1023),   
       .C_PROG_FULL_THRESH_ASSERT_VAL_WDCH (1023),   
       .C_PROG_FULL_THRESH_ASSERT_VAL_WRCH (1023),   
       .C_PROG_FULL_THRESH_ASSERT_VAL_RACH (1023),   
       .C_PROG_FULL_THRESH_ASSERT_VAL_RDCH (1023),   
       .C_PROG_FULL_THRESH_ASSERT_VAL_AXIS (1023),   
       .C_PROG_EMPTY_TYPE_WACH		(0),        
       .C_PROG_EMPTY_TYPE_WDCH		(0),        
       .C_PROG_EMPTY_TYPE_WRCH		(0),        
       .C_PROG_EMPTY_TYPE_RACH		(0),        
       .C_PROG_EMPTY_TYPE_RDCH		(0),        
       .C_PROG_EMPTY_TYPE_AXIS		(0),        
       .C_PROG_EMPTY_THRESH_ASSERT_VAL_WACH (1022),  
       .C_PROG_EMPTY_THRESH_ASSERT_VAL_WDCH (1022),  
       .C_PROG_EMPTY_THRESH_ASSERT_VAL_WRCH (1022),  
       .C_PROG_EMPTY_THRESH_ASSERT_VAL_RACH (1022),  
       .C_PROG_EMPTY_THRESH_ASSERT_VAL_RDCH (1022),  
       .C_PROG_EMPTY_THRESH_ASSERT_VAL_AXIS (1022),  
       .C_REG_SLICE_MODE_WACH		(0),        
       .C_REG_SLICE_MODE_WDCH		(0),        
       .C_REG_SLICE_MODE_WRCH		(0),        
       .C_REG_SLICE_MODE_RACH		(0),        
       .C_REG_SLICE_MODE_RDCH		(0),        
       .C_REG_SLICE_MODE_AXIS		(0)         
       )
     // }}} ---------------
     dist_ram_afifo_inst
      (.din                            (afifo_wdata),
       .rd_clk                         (phy_clk),
       .rd_en                          (afifo_rd),
       .rst                            (buf_phy_rst_q),
       .wr_clk                         (log_clk),
       .wr_en                          (afifo_wr),
       .almost_full                    (afifo_full),
       .dout                           (afifo_rdata),
       .empty                          (afifo_empty),
       .full                           (),
       .clk                            (),
       .int_clk                        (),
       .backup                         (),
       .backup_marker                  (),
       .prog_empty_thresh              (),
       .prog_empty_thresh_assert       (),
       .prog_empty_thresh_negate       (),
       .prog_full_thresh               (),
       .prog_full_thresh_assert        (),
       .prog_full_thresh_negate        (),
       .rd_rst                         (),
       .srst                           (),
       .wr_rst                         (),
       .almost_empty                   (),
       .data_count                     (),
       .overflow                       (),
       .prog_empty                     (),
       .prog_full                      (),
       .valid                          (),
       .rd_data_count                  (),
       .underflow                      (),
       .wr_ack                         (),
       .wr_data_count                  (),
       .sbiterr                        (),
       .dbiterr                        (),
       .injectsbiterr                  (),
       .injectdbiterr                  (),

       .sleep          (1'b0),// added with default values
       .wr_rst_busy    (),// added these 2 pins, core may not use those at the moment
       .rd_rst_busy    (),// added these 2 pins, core may not use those at the moment

       .m_aclk                         (),
       .s_aclk                         (),
       .s_aresetn                      (),
       .s_aclk_en                      (),
       .m_aclk_en                      (),
       .s_axi_awid                     (),
       .s_axi_awaddr                   (),
       .s_axi_awlen                    (),
       .s_axi_awsize                   (),
       .s_axi_awburst                  (),
       .s_axi_awlock                   (),
       .s_axi_awcache                  (),
       .s_axi_awprot                   (),
       .s_axi_awqos                    (),
       .s_axi_awregion                 (),
       .s_axi_awuser                   (),
       .s_axi_awvalid                  (),
       .s_axi_awready                  (),
       .s_axi_wid                      (),
       .s_axi_wdata                    (),
       .s_axi_wstrb                    (),
       .s_axi_wlast                    (),
       .s_axi_wuser                    (),
       .s_axi_wvalid                   (),
       .s_axi_wready                   (),
       .s_axi_bid                      (),
       .s_axi_bresp                    (),
       .s_axi_buser                    (),
       .s_axi_bvalid                   (),
       .s_axi_bready                   (),
       .m_axi_awid                     (),
       .m_axi_awaddr                   (),
       .m_axi_awlen                    (),
       .m_axi_awsize                   (),
       .m_axi_awburst                  (),
       .m_axi_awlock                   (),
       .m_axi_awcache                  (),
       .m_axi_awprot                   (),
       .m_axi_awqos                    (),
       .m_axi_awregion                 (),
       .m_axi_awuser                   (),
       .m_axi_awvalid                  (),
       .m_axi_awready                  (),
       .m_axi_wid                      (),
       .m_axi_wdata                    (),
       .m_axi_wstrb                    (),
       .m_axi_wlast                    (),
       .m_axi_wuser                    (),
       .m_axi_wvalid                   (),
       .m_axi_wready                   (),
       .m_axi_bid                      (),
       .m_axi_bresp                    (),
       .m_axi_buser                    (),
       .m_axi_bvalid                   (),
       .m_axi_bready                   (),
       .s_axi_arid                     (),
       .s_axi_araddr                   (),
       .s_axi_arlen                    (),
       .s_axi_arsize                   (),
       .s_axi_arburst                  (),
       .s_axi_arlock                   (),
       .s_axi_arcache                  (),
       .s_axi_arprot                   (),
       .s_axi_arqos                    (),
       .s_axi_arregion                 (),
       .s_axi_aruser                   (),
       .s_axi_arvalid                  (),
       .s_axi_arready                  (),
       .s_axi_rid                      (),
       .s_axi_rdata                    (),
       .s_axi_rresp                    (),
       .s_axi_rlast                    (),
       .s_axi_ruser                    (),
       .s_axi_rvalid                   (),
       .s_axi_rready                   (),
       .m_axi_arid                     (),
       .m_axi_araddr                   (),
       .m_axi_arlen                    (),
       .m_axi_arsize                   (),
       .m_axi_arburst                  (),
       .m_axi_arlock                   (),
       .m_axi_arcache                  (),
       .m_axi_arprot                   (),
       .m_axi_arqos                    (),
       .m_axi_arregion                 (),
       .m_axi_aruser                   (),
       .m_axi_arvalid                  (),
       .m_axi_arready                  (),
       .m_axi_rid                      (),
       .m_axi_rdata                    (),
       .m_axi_rresp                    (),
       .m_axi_rlast                    (),
       .m_axi_ruser                    (),
       .m_axi_rvalid                   (),
       .m_axi_rready                   (),
       .s_axis_tvalid                  (),
       .s_axis_tready                  (),
       .s_axis_tdata                   (),
       .s_axis_tstrb                   (),
       .s_axis_tkeep                   (),
       .s_axis_tlast                   (),
       .s_axis_tid                     (),
       .s_axis_tdest                   (),
       .s_axis_tuser                   (),
       .m_axis_tvalid                  (),
       .m_axis_tready                  (),
       .m_axis_tdata                   (),
       .m_axis_tstrb                   (),
       .m_axis_tkeep                   (),
       .m_axis_tlast                   (),
       .m_axis_tid                     (),
       .m_axis_tdest                   (),
       .m_axis_tuser                   (),
       .axi_aw_injectsbiterr           (),
       .axi_aw_injectdbiterr           (),
       .axi_aw_prog_full_thresh        (),
       .axi_aw_prog_empty_thresh       (),
       .axi_aw_data_count              (),
       .axi_aw_wr_data_count           (),
       .axi_aw_rd_data_count           (),
       .axi_aw_sbiterr                 (),
       .axi_aw_dbiterr                 (),
       .axi_aw_overflow                (),
       .axi_aw_underflow               (),
       .axi_aw_prog_full               (), // CR 724965 output port left with dummy assignment
       .axi_aw_prog_empty              (), // CR 724965 output port left with dummy assignment
       .axi_w_injectsbiterr            (),
       .axi_w_injectdbiterr            (),
       .axi_w_prog_full_thresh         (),
       .axi_w_prog_empty_thresh        (),
       .axi_w_data_count               (),
       .axi_w_wr_data_count            (),
       .axi_w_rd_data_count            (),
       .axi_w_sbiterr                  (),
       .axi_w_dbiterr                  (),
       .axi_w_overflow                 (),
       .axi_w_underflow                (),
       .axi_b_injectsbiterr            (),
       .axi_b_injectdbiterr            (),
       .axi_w_prog_full                (), // CR 724965 output port left with dummy assignment
       .axi_w_prog_empty               (), // CR 724965 output port left with dummy assignment
       .axi_b_prog_full_thresh         (),
       .axi_b_prog_empty_thresh        (),
       .axi_b_data_count               (),
       .axi_b_wr_data_count            (),
       .axi_b_rd_data_count            (),
       .axi_b_sbiterr                  (),
       .axi_b_dbiterr                  (),
       .axi_b_overflow                 (),
       .axi_b_underflow                (),
       .axi_ar_injectsbiterr           (),
       .axi_ar_injectdbiterr           (),
       .axi_b_prog_full                (), // CR 724965 output port left with dummy assignment
       .axi_b_prog_empty               (), // CR 724965 output port left with dummy assignment
       .axi_ar_prog_full_thresh        (),
       .axi_ar_prog_empty_thresh       (),
       .axi_ar_data_count              (),
       .axi_ar_wr_data_count           (),
       .axi_ar_rd_data_count           (),
       .axi_ar_sbiterr                 (),
       .axi_ar_dbiterr                 (),
       .axi_ar_overflow                (),
       .axi_ar_underflow               (),
       .axi_r_injectsbiterr            (),
       .axi_r_injectdbiterr            (),
       .axi_ar_prog_full               (),  // CR 724965 output port left with dummy assignment
       .axi_ar_prog_empty              (),  // CR 724965 output port left with dummy assignment
       .axi_r_prog_full_thresh         (),
       .axi_r_prog_empty_thresh        (),
       .axi_r_data_count               (),
       .axi_r_wr_data_count            (),
       .axi_r_rd_data_count            (),
       .axi_r_sbiterr                  (),
       .axi_r_dbiterr                  (),
       .axi_r_overflow                 (),
       .axi_r_underflow                (),
       .axis_injectsbiterr             (),
       .axis_injectdbiterr             (),
       .axi_r_prog_full                (),  // CR 724965 output port left with dummy assignment
       .axi_r_prog_empty               (),  // CR 724965 output port left with dummy assignment
       .axis_prog_full_thresh          (),
       .axis_prog_empty_thresh         (),
       .axis_data_count                (),
       .axis_wr_data_count             (),
       .axis_rd_data_count             (),
       .axis_sbiterr                   (),
       .axis_dbiterr                   (),
       .axis_overflow                  (),
       .axis_underflow                 (),
       .axis_prog_full                 (),  // CR 724965 output port left with dummy assignment
       .axis_prog_empty                ()   // CR 724965 output port left with dummy assignment
      );

    // }}} end Real Synch Unit ---
  end else                   begin: fake_sync_unit
    // {{{ Fake Synch Unit ---
    // in the case when no synchronization is required, simply connect the ins
    // to the outs.
    assign BTS_tx_data      = LD_buft_tdata;
    assign BTS_tx_start     = bts_buft_tstart;
    assign BTS_tx_last      = LD_buft_tlast;
    assign BTS_tx_valid     = LD_buft_tvalid;
    assign BTS_tx_keep      = {LD_buft_tkeep[5], LD_buft_tkeep[3], LD_buft_tkeep[1]};
    assign BTS_tx_user      = LD_buft_tuser;
    assign afifo_full       = 1'b0;

    always @ * begin
      BTS_buft_tready  = BT_tx_ready;
    end
    // }}} end Fake Synch Unit ---
  end
  endgenerate

  // {{{ Outstanding packets counter ---------

  // this piece of logic will be generated regardless of a unified clock or
  // not.  It keeps track of the total number of outstanding packets that have
  // been recieved by the buffer.  This is important to keep because we must
  // be able to reserve at least one final location for responses.

  // Synchronize the master enable signal before using.
  always @(posedge log_clk) begin
    if (buf_log_rst_q)
      pcfg_master_en_a <= #TCQ 1'b0;
    else
      pcfg_master_en_a <= #TCQ PC_master_enable;
  end

  // this is being done in order to prevent the tools from making two adders. This isn't as
  // easy to read but worth the cost savings. Add one when a new packet arrives. Subtract one
  // when the buffer logic sees an acknowledgement.
  assign outstanding_packets_inc = bts_buft_tstart && LD_buft_tvalid && BTS_buft_tready;
  assign outstanding_packets_dec = !log_packet_available_n;

  always @(posedge log_clk) begin
    if (buf_log_rst_q)
      BTS_response_only <= #TCQ 1'b0;
    // on an increment condition, evaluate for one less than the typical case
    else if (outstanding_packets_inc && !outstanding_packets_dec)
      BTS_response_only <= !pcfg_master_en_a ||
                             (outstanding_packets > (TX_DEPTH - RESPONSE_ONLY_THRESHOLD - 1));
    // typical case
    else
      BTS_response_only <= !pcfg_master_en_a ||
                             (outstanding_packets > (TX_DEPTH - RESPONSE_ONLY_THRESHOLD));
  end

  // either +1 or -1, depending on the operation
  wire [5:0] increment_value = outstanding_packets_inc ? 1 : -1;
  always @(posedge log_clk) begin
    if (buf_log_rst_q)
      outstanding_packets <= #TCQ 0;
    // if an incoming packet and an acknowledged packet arrive on the same cycle, they cancel out.
    else if (outstanding_packets_inc && !outstanding_packets_dec)
      outstanding_packets <= #TCQ outstanding_packets + increment_value; // +1 here
    else if (!outstanding_packets_inc && outstanding_packets_dec)
      outstanding_packets <= #TCQ outstanding_packets + increment_value; // -1 here
  end
  // }}} --------------------------------------


  // {{{ Start of Packet generation ----------

  always @(posedge log_clk) begin
    if (buf_log_rst_q)
      bts_buft_tstart <= #TCQ 1'b1;
    else if (LD_buft_tvalid && BTS_buft_tready)
      bts_buft_tstart <= #TCQ LD_buft_tlast;
  end
  // }}} --------------------------------------


  // {{{ Asynch FIFO for returning information from PHY domain --

  fifo_generator_vlog_beh
   // {{{ parameter list ---------------
   #(
     .C_COMMON_CLOCK                 (0),
     .C_COUNT_TYPE                   (0),
     .C_DATA_COUNT_WIDTH             (5),
     .C_DEFAULT_VALUE                ("BlankString"),
     .C_DIN_WIDTH                    (2),  // NOTE - CFR - this only needs to be 1
     .C_DOUT_RST_VAL                 ("0"),
     .C_DOUT_WIDTH                   (2),  // NOTE - CFR - this only needs to be 1
     .C_ENABLE_RLOCS                 (0),
     .C_ENABLE_RST_SYNC              (1),
     .C_ERROR_INJECTION_TYPE         (0),
     .C_FAMILY                       (C_FAMILY),
     .C_FULL_FLAGS_RST_VAL           (1),
     .C_HAS_ALMOST_EMPTY             (0),
     .C_HAS_ALMOST_FULL              (0),
     .C_HAS_BACKUP                   (0),
     .C_HAS_DATA_COUNT               (0),
     .C_HAS_INT_CLK                  (0),
     .C_HAS_MEMINIT_FILE             (0),
     .C_HAS_OVERFLOW                 (0),
     .C_HAS_RD_DATA_COUNT            (0),
     .C_HAS_RD_RST                   (0),
     .C_HAS_RST                      (1),
     .C_HAS_SRST                     (0),
     .C_HAS_UNDERFLOW                (0),
     .C_HAS_VALID                    (0),
     .C_HAS_WR_ACK                   (0),
     .C_HAS_WR_DATA_COUNT            (0),
     .C_HAS_WR_RST                   (0),
     .C_IMPLEMENTATION_TYPE          (2),
     .C_INIT_WR_PNTR_VAL             (0),
     .C_MEMORY_TYPE                  (2),
     .C_MIF_FILE_NAME                ("BlankString"),
     .C_MSGON_VAL                    (1),
     .C_OPTIMIZATION_MODE            (0),
     .C_OVERFLOW_LOW                 (0),
     .C_PRELOAD_LATENCY              (1),
     .C_PRELOAD_REGS                 (0),
     .C_PRIM_FIFO_TYPE               ("512x36"),
     .C_PROG_EMPTY_THRESH_ASSERT_VAL (2),
     .C_PROG_EMPTY_THRESH_NEGATE_VAL (3),
     .C_PROG_EMPTY_TYPE              (0),
     .C_PROG_FULL_THRESH_ASSERT_VAL  (29),
     .C_PROG_FULL_THRESH_NEGATE_VAL  (28),
     .C_PROG_FULL_TYPE               (0),
     .C_RD_DATA_COUNT_WIDTH          (5),
     .C_RD_DEPTH                     (TX_DEPTH),
     .C_RD_FREQ                      (1),
     .C_RD_PNTR_WIDTH                (PTR_WIDTH),
     .C_UNDERFLOW_LOW                (0),
     .C_USE_DOUT_RST                 (1),
     .C_USE_ECC                      (0),
     .C_USE_EMBEDDED_REG             (0),
     .C_USE_FIFO16_FLAGS             (0),
     .C_USE_FWFT_DATA_COUNT          (0),
     .C_VALID_LOW                    (0),
     .C_WR_ACK_LOW                   (0),
     .C_WR_DATA_COUNT_WIDTH          (5),
     .C_WR_DEPTH                     (TX_DEPTH),
     .C_WR_FREQ                      (1),
     .C_WR_PNTR_WIDTH                (PTR_WIDTH),
     .C_WR_RESPONSE_LATENCY          (1),
     
     //-- below parameters are newly added for v12_0, core doesnt use it
     //left @ default
     .C_USE_PIPELINE_REG	(0),		// --
     .C_POWER_SAVING_MODE	(0),		// --
     .C_SYNCHRONIZER_STAGE	(2),		// --
     .C_INTERFACE_TYPE	(0),		// --
     .C_AXI_TYPE		(1),		// --
     .C_HAS_AXI_WR_CHANNEL	(1),		// --
     .C_HAS_AXI_RD_CHANNEL	(1),		// --
     .C_HAS_SLAVE_CE		(0),		// --
     .C_HAS_MASTER_CE		(0),		// --
     .C_ADD_NGC_CONSTRAINT	(0),		// --
     .C_USE_COMMON_OVERFLOW	(0),		// --
     .C_USE_COMMON_UNDERFLOW	(0),		// --
     .C_USE_DEFAULT_SETTINGS	(0),		// --
     .C_AXI_ID_WIDTH		(1),		// --
     .C_AXI_ADDR_WIDTH	(32),		// --
     .C_AXI_DATA_WIDTH	(64),		// --
     .C_AXI_LEN_WIDTH		(8),		// --
     .C_AXI_LOCK_WIDTH	(1),		// --
     .C_HAS_AXI_ID		(0),		// --
     .C_HAS_AXI_AWUSER	(0),		// --
     .C_HAS_AXI_WUSER		(0),		// --
     .C_HAS_AXI_BUSER		(0),		// --
     .C_HAS_AXI_ARUSER	(0),		// --
     .C_HAS_AXI_RUSER		(0),		// --
     .C_AXI_ARUSER_WIDTH	(1),		// --
     .C_AXI_AWUSER_WIDTH	(1),		// --
     .C_AXI_WUSER_WIDTH	(1),		// --
     .C_AXI_BUSER_WIDTH	(1),		// --
     .C_AXI_RUSER_WIDTH	(1),		// --
     .C_HAS_AXIS_TDATA	(1),		// --
     .C_HAS_AXIS_TID		(0),		// --
     .C_HAS_AXIS_TDEST	(0),		// --
     .C_HAS_AXIS_TUSER	(1),		// --
     .C_HAS_AXIS_TREADY	(1),		// --
     .C_HAS_AXIS_TLAST	(0),		// --
     .C_HAS_AXIS_TSTRB	(0),		// --
     .C_HAS_AXIS_TKEEP	(0),		// --
     .C_AXIS_TDATA_WIDTH	(8),		// --
     .C_AXIS_TID_WIDTH	(1),		// --
     .C_AXIS_TDEST_WIDTH	(1),		// --
     .C_AXIS_TUSER_WIDTH	(4),		// --
     .C_AXIS_TSTRB_WIDTH	(1),		// --
     .C_AXIS_TKEEP_WIDTH	(1),		// --
     .C_WACH_TYPE		(0),		// --
     .C_WDCH_TYPE		(0),		// --
     .C_WRCH_TYPE		(0),		// --
     .C_RACH_TYPE		(0),		// --
     .C_RDCH_TYPE		(0),		// --
     .C_AXIS_TYPE		(0),		// --
     .C_IMPLEMENTATION_TYPE_WACH (1),	// --
     .C_IMPLEMENTATION_TYPE_WDCH (1),	// --
     .C_IMPLEMENTATION_TYPE_WRCH (1),	// --
     .C_IMPLEMENTATION_TYPE_RACH (1),	// --
     .C_IMPLEMENTATION_TYPE_RDCH (1),	// --
     .C_IMPLEMENTATION_TYPE_AXIS (1),	// --
     .C_APPLICATION_TYPE_WACH	(0),	// --
     .C_APPLICATION_TYPE_WDCH	(0),	// --
     .C_APPLICATION_TYPE_WRCH	(0),	// --
     .C_APPLICATION_TYPE_RACH	(0),	// --
     .C_APPLICATION_TYPE_RDCH	(0),	// --
     .C_APPLICATION_TYPE_AXIS	(0),	// --
     .C_PRIM_FIFO_TYPE_WACH	("512x36"),	// --
     .C_PRIM_FIFO_TYPE_WDCH	("1kx36"),	// --
     .C_PRIM_FIFO_TYPE_WRCH	("512x36"),	// --
     .C_PRIM_FIFO_TYPE_RACH	("512x36"),	// --
     .C_PRIM_FIFO_TYPE_RDCH	("1kx36"),	// --
     .C_PRIM_FIFO_TYPE_AXIS	("1kx18"),	// --
     .C_USE_ECC_WACH		(0),		// --
     .C_USE_ECC_WDCH		(0),		// --
     .C_USE_ECC_WRCH		(0),		// --
     .C_USE_ECC_RACH		(0),		// --
     .C_USE_ECC_RDCH		(0),		// --
     .C_USE_ECC_AXIS		(0),		// --
     .C_ERROR_INJECTION_TYPE_WACH (0),	// --
     .C_ERROR_INJECTION_TYPE_WDCH (0),	// --
     .C_ERROR_INJECTION_TYPE_WRCH (0),	// --
     .C_ERROR_INJECTION_TYPE_RACH (0),	// --
     .C_ERROR_INJECTION_TYPE_RDCH (0),	// --
     .C_ERROR_INJECTION_TYPE_AXIS (0),	// --
     .C_DIN_WIDTH_WACH	(32),		// --
     .C_DIN_WIDTH_WDCH	(64),		// --
     .C_DIN_WIDTH_WRCH	(2),		// --
     .C_DIN_WIDTH_RACH	(32),		// --
     .C_DIN_WIDTH_RDCH	(64),		// --
     .C_DIN_WIDTH_AXIS	(1),		// --
     .C_WR_DEPTH_WACH		(16),		// --
     .C_WR_DEPTH_WDCH		(1024),		// --
     .C_WR_DEPTH_WRCH		(16),		// --
     .C_WR_DEPTH_RACH		(16),		// --
     .C_WR_DEPTH_RDCH		(1024),		// --
     .C_WR_DEPTH_AXIS		(1024),		// --
     .C_WR_PNTR_WIDTH_WACH	(4),	// --
     .C_WR_PNTR_WIDTH_WDCH	(10),	// --
     .C_WR_PNTR_WIDTH_WRCH	(4),	// --
     .C_WR_PNTR_WIDTH_RACH	(4),	// --
     .C_WR_PNTR_WIDTH_RDCH	(10),	// --
     .C_WR_PNTR_WIDTH_AXIS	(10),	// --
     .C_HAS_DATA_COUNTS_WACH	(0),	// --
     .C_HAS_DATA_COUNTS_WDCH	(0),	// --
     .C_HAS_DATA_COUNTS_WRCH	(0),	// --
     .C_HAS_DATA_COUNTS_RACH	(0),	// --
     .C_HAS_DATA_COUNTS_RDCH	(0),	// --
     .C_HAS_DATA_COUNTS_AXIS	(0),	// --
     .C_HAS_PROG_FLAGS_WACH	(0),	// --
     .C_HAS_PROG_FLAGS_WDCH	(0),	// --
     .C_HAS_PROG_FLAGS_WRCH	(0),	// --
     .C_HAS_PROG_FLAGS_RACH	(0),	// --
     .C_HAS_PROG_FLAGS_RDCH	(0),	// --
     .C_HAS_PROG_FLAGS_AXIS	(0),	// --
     .C_PROG_FULL_TYPE_WACH	(0),	// --
     .C_PROG_FULL_TYPE_WDCH	(0),	// --
     .C_PROG_FULL_TYPE_WRCH	(0),	// --
     .C_PROG_FULL_TYPE_RACH	(0),	// --
     .C_PROG_FULL_TYPE_RDCH	(0),	// --
     .C_PROG_FULL_TYPE_AXIS	(0),	// --
     .C_PROG_FULL_THRESH_ASSERT_VAL_WACH (1023),// --
     .C_PROG_FULL_THRESH_ASSERT_VAL_WDCH (1023),// --
     .C_PROG_FULL_THRESH_ASSERT_VAL_WRCH (1023),// --
     .C_PROG_FULL_THRESH_ASSERT_VAL_RACH (1023),// --
     .C_PROG_FULL_THRESH_ASSERT_VAL_RDCH (1023),// --
     .C_PROG_FULL_THRESH_ASSERT_VAL_AXIS (1023),// --
     .C_PROG_EMPTY_TYPE_WACH	(0),	// --
     .C_PROG_EMPTY_TYPE_WDCH	(0),	// --
     .C_PROG_EMPTY_TYPE_WRCH	(0),	// --
     .C_PROG_EMPTY_TYPE_RACH	(0),	// --
     .C_PROG_EMPTY_TYPE_RDCH	(0),	// --
     .C_PROG_EMPTY_TYPE_AXIS	(0),	// --
     .C_PROG_EMPTY_THRESH_ASSERT_VAL_WACH (1022),// --
     .C_PROG_EMPTY_THRESH_ASSERT_VAL_WDCH (1022),// --
     .C_PROG_EMPTY_THRESH_ASSERT_VAL_WRCH (1022),// --
     .C_PROG_EMPTY_THRESH_ASSERT_VAL_RACH (1022),// --
     .C_PROG_EMPTY_THRESH_ASSERT_VAL_RDCH (1022),// --
     .C_PROG_EMPTY_THRESH_ASSERT_VAL_AXIS (1022),// --
     .C_REG_SLICE_MODE_WACH	(0),	// --
     .C_REG_SLICE_MODE_WDCH	(0),	// --
     .C_REG_SLICE_MODE_WRCH	(0),	// --
     .C_REG_SLICE_MODE_RACH	(0),	// --
     .C_REG_SLICE_MODE_RDCH	(0),	// --
     .C_REG_SLICE_MODE_AXIS	(0)	// --
     )
   // }}} ---------------
   srl16_fifo_inst
      (/*.din                            (2'b1),  // NOTE - CFR - This only needs to be 1
       .rd_clk                         (log_clk),
       .rd_en                          (outstanding_packets_dec),
       .rst                            (buf_phy_rst_q),
       .wr_clk                         (phy_clk),
       .wr_en                          (BT_packet_ack),
       .dout                           (),
       .empty                          (log_packet_available_n),
      */
        .backup                         (),
        .backup_marker                  (),
        .clk                            (),
        .rst                            (buf_phy_rst_q),
        .srst                           (),
        .wr_clk                         (phy_clk),
        .wr_rst                         (),
        .rd_clk                         (log_clk),
        .rd_rst                         (),
        .din                            (2'b1),
        .wr_en                          (BT_packet_ack),
        .rd_en                          (outstanding_packets_dec),
        .prog_empty_thresh              (),
        .prog_empty_thresh_assert       (),
        .prog_empty_thresh_negate       (),
        .prog_full_thresh               (),
        .prog_full_thresh_assert        (),
        .prog_full_thresh_negate        (),
        .int_clk                        (),
        .injectdbiterr                  (),
        .injectsbiterr                  (),
        .sleep                          (1'b0),
        .dout                           (),
        .full                           (),
        .almost_full                    (),
        .wr_ack                         (),
        .overflow                       (),
        .empty                          (log_packet_available_n),
        .almost_empty                   (),
        .valid                          (),
        .underflow                      (),
        .data_count                     (),
        .rd_data_count                  (),
        .wr_data_count                  (),
        .prog_full                      (),
        .prog_empty                     (),
        .sbiterr                        (),
        .dbiterr                        (),
        .wr_rst_busy                    (),
        .rd_rst_busy                    (),
        .m_aclk                         (),
        .s_aclk                         (),
        .s_aresetn                      (),
        .s_aclk_en                      (),
        .m_aclk_en                      (),
        
        .s_axi_awid                     (),
        .s_axi_awaddr                   (),
        .s_axi_awlen                    (),
        .s_axi_awsize                   (),
        .s_axi_awburst                  (),
        .s_axi_awlock                   (),
        .s_axi_awcache                  (),
        .s_axi_awprot                   (),
        .s_axi_awqos                    (),
        .s_axi_awregion                 (),
        .s_axi_awuser                   (),
        .s_axi_awvalid                  (),
        .s_axi_awready                  (),
        .s_axi_wid                      (),
        .s_axi_wdata                    (),
        .s_axi_wstrb                    (),
        .s_axi_wlast                    (),
        .s_axi_wuser                    (),
        .s_axi_wvalid                   (),
        .s_axi_wready                   (),
        .s_axi_bid                      (),
        .s_axi_bresp                    (),
        .s_axi_buser                    (),
        .s_axi_bvalid                   (),
        .s_axi_bready                   (),
        
        .m_axi_awid                     (),
        .m_axi_awaddr                   (),
        .m_axi_awlen                    (),
        .m_axi_awsize                   (),
        .m_axi_awburst                  (),
        .m_axi_awlock                   (),
        .m_axi_awcache                  (),
        .m_axi_awprot                   (),
        .m_axi_awqos                    (),
        .m_axi_awregion                 (),
        .m_axi_awuser                   (),
        .m_axi_awvalid                  (),
        .m_axi_awready                  (),
        .m_axi_wid                      (),
        .m_axi_wdata                    (),
        .m_axi_wstrb                    (),
        .m_axi_wlast                    (),
        .m_axi_wuser                    (),
        .m_axi_wvalid                   (),
        .m_axi_wready                   (),
        .m_axi_bid                      (),
        .m_axi_bresp                    (),
        .m_axi_buser                    (),
        .m_axi_bvalid                   (),
        .m_axi_bready                   (),
        
        .s_axi_arid                     (),
        .s_axi_araddr                   (), 
        .s_axi_arlen                    (),
        .s_axi_arsize                   (),
        .s_axi_arburst                  (),
        .s_axi_arlock                   (),
        .s_axi_arcache                  (),
        .s_axi_arprot                   (),
        .s_axi_arqos                    (),
        .s_axi_arregion                 (),
        .s_axi_aruser                   (),
        .s_axi_arvalid                  (),
        .s_axi_arready                  (),
        .s_axi_rid                      (),       
        .s_axi_rdata                    (), 
        .s_axi_rresp                    (),
        .s_axi_rlast                    (),
        .s_axi_ruser                    (),
        .s_axi_rvalid                   (),
        .s_axi_rready                   (),
        
        .m_axi_arid                     (),        
        .m_axi_araddr                   (),  
        .m_axi_arlen                    (),
        .m_axi_arsize                   (),
        .m_axi_arburst                  (),
        .m_axi_arlock                   (),
        .m_axi_arcache                  (),
        .m_axi_arprot                   (),
        .m_axi_arqos                    (),
        .m_axi_arregion                 (),
        .m_axi_aruser                   (),
        .m_axi_arvalid                  (),
        .m_axi_arready                  (),
        .m_axi_rid                      (),        
        .m_axi_rdata                    (),  
        .m_axi_rresp                    (),
        .m_axi_rlast                    (),
        .m_axi_ruser                    (),
        .m_axi_rvalid                   (),
        .m_axi_rready                   (),
        
        .s_axis_tvalid                  (),
        .s_axis_tready                  (),
        .s_axis_tdata                   (),
        .s_axis_tstrb                   (),
        .s_axis_tkeep                   (),
        .s_axis_tlast                   (),
        .s_axis_tid                     (),
        .s_axis_tdest                   (),
        .s_axis_tuser                   (),
        
        .m_axis_tvalid                  (),
        .m_axis_tready                  (),
        .m_axis_tdata                   (),
        .m_axis_tstrb                   (),
        .m_axis_tkeep                   (),
        .m_axis_tlast                   (),
        .m_axis_tid                     (),
        .m_axis_tdest                   (),
        .m_axis_tuser                   (),
        
        .axi_aw_injectsbiterr           (),
        .axi_aw_injectdbiterr           (),
        .axi_aw_prog_full_thresh        (),
        .axi_aw_prog_empty_thresh       (),
        .axi_aw_data_count              (),
        .axi_aw_wr_data_count           (),
        .axi_aw_rd_data_count           (),
        .axi_aw_sbiterr                 (),
        .axi_aw_dbiterr                 (),
        .axi_aw_overflow                (),
        .axi_aw_underflow               (),
        .axi_aw_prog_full               (),
        .axi_aw_prog_empty              (),
        
        .axi_w_injectsbiterr            (),
        .axi_w_injectdbiterr            (),
        .axi_w_prog_full_thresh         (),
        .axi_w_prog_empty_thresh        (),
        .axi_w_data_count               (),
        .axi_w_wr_data_count            (),
        .axi_w_rd_data_count            (),
        .axi_w_sbiterr                  (),
        .axi_w_dbiterr                  (),
        .axi_w_overflow                 (),
        .axi_w_underflow                (),
        .axi_w_prog_full                (),
        .axi_w_prog_empty               (),
        
        .axi_b_injectsbiterr            (),
        .axi_b_injectdbiterr            (),
        .axi_b_prog_full_thresh         (),
        .axi_b_prog_empty_thresh        (),
        .axi_b_data_count               (),
        .axi_b_wr_data_count            (),
        .axi_b_rd_data_count            (),
        .axi_b_sbiterr                  (),
        .axi_b_dbiterr                  (),
        .axi_b_overflow                 (),
        .axi_b_underflow                (),
        .axi_b_prog_full                (),
        .axi_b_prog_empty               (),
        
        .axi_ar_injectsbiterr           (),
        .axi_ar_injectdbiterr           (),
        .axi_ar_prog_full_thresh        (),
        .axi_ar_prog_empty_thresh       (),
        .axi_ar_data_count              (),
        .axi_ar_wr_data_count           (),
        .axi_ar_rd_data_count           (),
        .axi_ar_sbiterr                 (),
        .axi_ar_dbiterr                 (),
        .axi_ar_overflow                (),
        .axi_ar_underflow               (),
        .axi_ar_prog_full               (),
        .axi_ar_prog_empty              (),
        
        .axi_r_injectsbiterr            (),
        .axi_r_injectdbiterr            (),
        .axi_r_prog_full_thresh         (),
        .axi_r_prog_empty_thresh        (),
        .axi_r_data_count               (),
        .axi_r_wr_data_count            (),
        .axi_r_rd_data_count            (),
        .axi_r_sbiterr                  (),
        .axi_r_dbiterr                  (),
        .axi_r_overflow                 (),
        .axi_r_underflow                (),
        .axi_r_prog_full                (),
        .axi_r_prog_empty               (),
        
        .axis_injectsbiterr             (),
        .axis_injectdbiterr             (),
        .axis_prog_full_thresh          (),
        .axis_prog_empty_thresh         (),
        .axis_data_count                (),
        .axis_wr_data_count             (),
        .axis_rd_data_count             (),
        .axis_sbiterr                   (),
        .axis_dbiterr                   (),
        .axis_overflow                  (),
        .axis_underflow                 (),
        .axis_prog_full                 (),
        .axis_prog_empty                ()

  );

  // }}} -----------------------------------

endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/buf/srio_gen2_v4_1_16_buf_tx_bram_bank.v#1 $
//
// BUF_TX_BRAM_BANK
// Description:
// This module instantiates a family-specific memory module. It calls
// BLK_MEM_GEN from Coregen
//
// Hierarchy:
// BUF_TOP
//  |______BUF_TX
//  |____________BUF_TX_SYNC_UNIT
//  |____________BUF_TX_BRAM_BANK <-- this module
//  |______BUF_RX
//  |____________BUF_RX_ASYNC_PASSAGE
//  |____________BUF_RX_BRAM_BANK
//----------------------------------------------------------------------
`timescale 1ps/1ps
(* DowngradeIPIdentifiedWarnings = "yes" *)

module srio_gen2_v4_1_16_buf_tx_bram_bank
  #(
    parameter TCQ           = 100,
    parameter C_FAMILY      = "virtex6",         // {virtex5, virtex6, virtex7, spartan6, spartan7}
    parameter C_INDEX_LEN   = 6,                 // {6}
    parameter C_ADDR_LEN    = 11)                // {9, 10, 11}
   (
   // {{{ port declarations -----------------
    input                   phy_clk,             // Physical Layer clock
    input                   buf_phy_rst_q,       // Synchronous Phy Layer reset
    // in from tx buffer
    input [C_ADDR_LEN-1:0]  BT_bram_waddr,       // Write address for memory
    input                   BT_bram_rd,          // Read enable
    input [C_ADDR_LEN-1:0]  BT_bram_raddr,       // Read address for memory
    input                   BT_bram_we,          // Write enable
    // in from synchronization unit
    input [63:0]            BTS_tx_data,         // Data In
    input  [1:0]            BTS_tx_user,         // User Field
    input                   BTS_tx_start,        // Start of Frame
    input                   BTS_tx_last,         // End of Frame
    input  [2:0]            BTS_tx_keep,         // Remainder
    // out to Physical layer
    output [63:0]           BTB_tx_bram_data,    // Data Out
    output [1:0]            BTB_tx_bram_user,    // User Field
    output                  BTB_tx_bram_start,   // Start of Frame
    output                  BTB_tx_bram_last,    // End of Frame
    output [2:0]            BTB_tx_bram_keep     // Remainder
   // }}} ---------------------------------
   );


  // {{{ local parameters ------------------
  localparam C_MEM_DEPTH = 1 << C_ADDR_LEN;
  // }}} ---------------------------------


  // {{{ wire declarations -----------------
  wire [70:0] bram_data_in  = {BTS_tx_keep, BTS_tx_last, BTS_tx_start, BTS_tx_user, BTS_tx_data};
  wire [70:0] bram_data_out;

  assign {BTB_tx_bram_keep, BTB_tx_bram_last, BTB_tx_bram_start, BTB_tx_bram_user, BTB_tx_bram_data}  = bram_data_out;

    // *- COVERAGE (BT_mask_false_last)
    // observe a false last being masked

  // }}} ---------------------------------


  // {{{ Block memory Instantiation --------
  blk_mem_gen_v8_4_4                                          // blk_mem_gen_v8_0 values
   #(
     .C_ADDRA_WIDTH                 (C_ADDR_LEN),           // (C_ADDR_LEN),          
     .C_ADDRB_WIDTH                 (C_ADDR_LEN),           // (C_ADDR_LEN),          
     .C_ALGORITHM                   (1),                    // (1),                   
     .C_AXI_ID_WIDTH                (4),                    // (4),                   
     .C_AXI_SLAVE_TYPE              (4),                    // (4),                   
     .C_AXI_TYPE                    (4),                    // (4),                   
     .C_BYTE_SIZE                   (9),                    // (9),                   
     .C_COMMON_CLK                  (1),                    // (1),                   
     .C_DEFAULT_DATA                ("0"),                  // ("0"),                 
     .C_DISABLE_WARN_BHV_COLL       (0),                    // (0),                   
     .C_DISABLE_WARN_BHV_RANGE      (1),                    // (1),                   
     .C_ELABORATION_DIR             (""),                   // (""),                  
     .C_ENABLE_32BIT_ADDRESS        (0),                    // (0),                   
     .C_FAMILY                      (C_FAMILY),             // (C_FAMILY),            

     .C_HAS_AXI_ID                  (0),                    // not present in this instance 

     .C_HAS_ENA                     (1),                    // (1),                   
     .C_HAS_ENB                     (1),                    // (1),                   
     .C_HAS_INJECTERR               (0),                    // (0),                   
     .C_HAS_MEM_OUTPUT_REGS_A       (0),                    // (0),                   
     .C_HAS_MEM_OUTPUT_REGS_B       (0),                    // (0),                   
     .C_HAS_MUX_OUTPUT_REGS_A       (0),                    // (0),                   
     .C_HAS_MUX_OUTPUT_REGS_B       (0),                    // (0),                   
     .C_HAS_REGCEA                  (0),                    // (0),                   
     .C_HAS_REGCEB                  (0),                    // (0),                   
     .C_HAS_RSTA                    (0),                    // (0),                   
     .C_HAS_RSTB                    (1),                    // (1),                   
     .C_HAS_SOFTECC_INPUT_REGS_A    (0),                    // (0),                   
     .C_HAS_SOFTECC_OUTPUT_REGS_B   (0),                    // (0),                   
     .C_INITA_VAL                   ("0"),                  // ("0"),                 
     .C_INITB_VAL                   ("0"),                  // ("0"),                 
     .C_INTERFACE_TYPE              (0),                    // (0),                   
     .C_INIT_FILE_NAME              ("no_coe_file_loaded"), // ("no_coe_file_loaded"),
     .C_LOAD_INIT_FILE              (0),                    // (0),                   
     .C_MEM_TYPE                    (1),                    // (1),                   
     .C_MUX_PIPELINE_STAGES         (0),                    // (0),                   
     .C_PRIM_TYPE                   (1),                    // (1),                   
     .C_READ_DEPTH_A                (C_MEM_DEPTH),          // (C_MEM_DEPTH),         
     .C_READ_DEPTH_B                (C_MEM_DEPTH),          // (C_MEM_DEPTH),         
     .C_READ_WIDTH_A                (71),                   // (71),                  
     .C_READ_WIDTH_B                (71),                   // (71),                  
     .C_RSTRAM_A                    (0),                    // (0),                   
     .C_RSTRAM_B                    (0),                    // (0),                   
     .C_RST_PRIORITY_A              ("CE"),                 // ("CE"),                
     .C_RST_PRIORITY_B              ("CE"),                 // ("CE"),                
     //.C_RST_TYPE                    ("SYNC"),               // ("SYNC"),-- assigned default value in the fifo_generator_v12_0 core              
     .C_SIM_COLLISION_CHECK         ("ALL"),                // ("ALL"),               
     .C_USE_BYTE_WEA                (0),                    // (0),                   
     .C_USE_BYTE_WEB                (0),                    // (0),                   
     .C_USE_DEFAULT_DATA            (0),                    // (0),                   
     .C_USE_ECC                     (0),                    // (0),                   
     .C_USE_SOFTECC                 (0),                    // (0),                   
     .C_WEA_WIDTH                   (1),                    // (1),                   
     .C_WEB_WIDTH                   (1),                    // (1),                   
     .C_WRITE_DEPTH_A               (C_MEM_DEPTH),          // (C_MEM_DEPTH),         
     .C_WRITE_DEPTH_B               (C_MEM_DEPTH),          // (C_MEM_DEPTH),         
     .C_WRITE_MODE_A                ("WRITE_FIRST"),        // ("WRITE_FIRST"),       
     .C_WRITE_MODE_B                ("WRITE_FIRST"),        // ("WRITE_FIRST"),       
     .C_WRITE_WIDTH_A               (71),                   // (71),                  
     .C_WRITE_WIDTH_B               (71),                   // (71),                  
     .C_XDEVICEFAMILY               (C_FAMILY),             // (C_FAMILY))

     // newly added parameters for the Diablo/US updates, leave default // 1/13/2015
     .C_USE_URAM                    (0),
     .C_EN_SAFETY_CKT               (0),
     .C_EN_DEEPSLEEP_PIN	    (0),
     .C_EN_SHUTDOWN_PIN	            (0),
     .C_EN_RDADDRA_CHG	            (0),
     .C_EN_RDADDRB_CHG	            (0)


     //_____________Below are newly added with blk_mem_gen_v8_2 version
     //_____________as per block mem gen owner, can be left at default or
     //_____________not included in the instance
     // .C_USE_BRAM_BLOCK		(0),
     // .C_CTRL_ECC_ALGO		("NONE"),
     // .C_INIT_FILE		("blk_mem_gen_0.mem"),
     // .C_EN_ECC_PIPE		(0),
     // .C_EN_SLEEP_PIN		(0),
     // .C_COUNT_36K_BRAM		("0"),
     // .C_COUNT_18K_BRAM		("1"),
     // .C_EST_POWER_SUMMARY	("Estimated Power for IP     :     3.0361 mW")
     )                                                       
   blk_mem_inst
    (
     .clka                        (phy_clk),
     .dina                        (bram_data_in),
     .addra                       (BT_bram_waddr),
     .ena                         (1'b1),
     .regcea                      (1'b0),
     .wea                         (BT_bram_we),
     .rsta                        (buf_phy_rst_q),
     .douta                       (),
     .clkb                        (phy_clk),
     .dinb                        (71'h0),
     .addrb                       (BT_bram_raddr),
     .enb                         (BT_bram_rd),
     .regceb                      (1'b0),
     .web                         (1'b0),
     .rstb                        (buf_phy_rst_q),
     .doutb                       (bram_data_out),
     .sbiterr                     (),
     .dbiterr                     (),
     .injectsbiterr               (),
     .injectdbiterr               (),
     .rdaddrecc                   (),

   // dont touch ports, new addition with default drive, // 1/13/2015
     .deepsleep                   (1'b0),
     .shutdown                    (1'b0),

     .s_aclk                      (),
     .s_aresetn                   (),
     .s_axi_awid                  (),
     .s_axi_awaddr                (),
     .s_axi_awlen                 (),
     .s_axi_awsize                (),
     .s_axi_awburst               (),
     .s_axi_awvalid               (),
     .s_axi_awready               (),
     .s_axi_wdata                 (),
     .s_axi_wstrb                 (),
     .s_axi_wlast                 (),
     .s_axi_wvalid                (),
     .s_axi_wready                (),
     .s_axi_bid                   (),
     .s_axi_bresp                 (),
     .s_axi_bvalid                (),
     .s_axi_bready                (),
     .s_axi_arid                  (),
     .s_axi_araddr                (),
     .s_axi_arlen                 (),
     .s_axi_arsize                (),
     .s_axi_arburst               (),
     .s_axi_arvalid               (),
     .s_axi_arready               (),
     .s_axi_rid                   (),
     .s_axi_rdata                 (),
     .s_axi_rresp                 (),
     .s_axi_rlast                 (),
     .s_axi_rvalid                (),
     .s_axi_rready                (),
     .s_axi_injectsbiterr         (),
     .s_axi_injectdbiterr         (),
     .s_axi_sbiterr               (),
     .s_axi_dbiterr               (),
     .s_axi_rdaddrecc               (),
     .sleep                       (1'b0),
     .eccpipece                   (1'b0)

    );
    
  // }}} ---------------------------------


endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//---------------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/log/srio_gen2_v4_1_16_log_top.v#1 $
//---------------------------------------------------------------------------
`timescale 1ps/1ps
// ------------------------------------------------
// below attribute is added to supress the synthesis warnings in vivado tool 8:3332
(* DowngradeIPIdentifiedWarnings="yes" *)
// ------------------------------------------------


module srio_gen2_v4_1_16_log_top #(
  // {{{ LOG Parameters
  parameter TCQ                       = 100,         // in ps
  parameter EVAL                      = 1,           // Includes the evaluation timer
  parameter DEVICEID_WIDTH            = 8,           // Indicates Source/Dest ID width {8, 16}
  parameter DEVICEID                  = 16'h00FF,    // Reset value for the DeviceID register {16'h0 - 16'hFFFF}
  parameter INIT_NREAD                = 1,           // If 1, core may initiate NRead transactions {0, 1}
  parameter INIT_NWRITE               = 1,           // If 1, core may initiate NWrite transactions {0, 1}
  parameter INIT_NWRITE_R             = 1,           // If 1, core may initiate NWrite_R transactions {0, 1}
  parameter INIT_SWRITE               = 1,           // If 1, core may initiate SWrite transactions {0, 1}
  parameter INIT_DB                   = 1,           // If 1, core may initiate Doorbell transactions {0, 1}
  parameter INIT_DS                   = 1,           // If 1, core may initiate Data Streaming {0, 1}
  parameter INIT_ATOMIC               = 1,           // If 1, core may initiate Atomic transactions {0, 1}
  parameter TARGET_NREAD              = 1,           // If 1, core may sink NRead transactions {0, 1}
  parameter TARGET_NWRITE             = 1,           // If 1, core may sink NWrite transactions {0, 1}
  parameter TARGET_NWRITE_R           = 1,           // If 1, core may sink NWrite_R transactions {0, 1}
  parameter TARGET_SWRITE             = 1,           // If 1, core may sink SWrite transactions {0, 1}
  parameter TARGET_DB                 = 1,           // If 1, core may sink Doorbell transactions {0, 1}
  parameter TARGET_DS                 = 1,           // If 1, core may sink Data Streaming {0, 1}
  parameter TARGET_ATOMIC             = 1,           // If 1, core may sink Atomic transactions {0, 1}
  parameter MSG_INIT_SINGLE           = 1,           // If 1, core may initiate single segment msg transactions {0, 1}
  parameter MSG_INIT_MULTI            = 1,           // If 1, core may initiate multi-segment msg transactions {0, 1}
  parameter MSG_SINK_SINGLE           = 1,           // If 1, core may sink single segment msg transactions {0, 1}
  parameter MSG_SINK_MULTI            = 1,           // If 1, core may sink multi-segment msg transactions {0, 1}
  parameter CRF_SUPPORT               = 1,           // If set, the core supports use of the CRF flag {0,1}
  parameter SINGLE_SEG_MBOX           = 16,          // Number of single segment mailboxes to support {0 - 64}
  parameter MAINT_SOURCE              = 1,           // If 1, core may source maint transactions {0, 1}
  parameter MAINT_CFG                 = 1,           // If 1, log maint block exists {0, 1}
  parameter DEVID_CAR                 = 32'h00000000,// Reset value for Device Identity CAR {32�h00000000�?32�hFFFFFFFF}
  parameter DEVINFO_CAR               = 32'h00000000,// Reset value for Device Info CAR {32�h00000000�?32�hFFFFFFFF}
  parameter DEV_CAR_OVRD              = 0,           // If 1, DEV*CAR param values used {0,1}
  parameter LCSBA_SUPPORT             = 1,           // If 1, indicates the LCSBA is used {0, 1}
  parameter LCSBA                     = 10'h3FF,     // Reset value for LCSBA register {0 - 10'h3FF}
  parameter HW_ARCH                   = 2,           // Device {V5LXT(0), V5FXT(1), V6LXT(2), V6CXT(3), S6LXT(4)}
  parameter ASSY_ID                   = 16'h0,       // Assembly ID from GUI {16'h0 - 16'hFFFF}
  parameter ASSY_VENDOR               = 16'h0,       // Assembly Vendor ID  {16'h0 - 16'hFFFF}
  parameter ASSY_REV                  = 16'h0,       // Assembly Revision {16'h0 - 16'hFFFF}
  parameter PHY_EF_PTR                = 16'h0100,    // Extended Features pointer {16'h0 - 16'hFFFF}
  parameter PE_BRIDGE                 = 0,           // PE is a bridge {0, 1}
  parameter PE_MEMORY                 = 1,           // PE is a memory {0, 1}
  parameter PE_PROC                   = 0,           // PE is a processor {0, 1}
  parameter PE_SWITCH                 = 0,           // PE is a switch {0, 1}
  parameter VC                        = 0,           // VC Support {0, 1}
  parameter PORT_IO_HELLO             = 1,           // The I/O ports use HELLO format {0,1}
  parameter PORT_MSG_HELLO            = 1,           // The Messaging ports use HELLO format {0,1}
  parameter PORT_MAINT_HELLO          = 1,           // The Maintenance ports use HELLO format {0,1}
  parameter PORT_IO_STYLE             = 1,           // 0: Condensed I/O style; 1: Init/Targ style; 2: Rd/Wr {0-2}
  parameter PORT_MSG_STYLE            = 1,           // MSGs go to 0: I/O port (msg ports disabled);
                                                       //            1: MSG port; 2: UserDef {0-2}
  parameter PORT_MAINT_STYLE          = 1,           // MAINTs go to 0: I/O port (maint ports disabled);
                                                       //              1: MAINT port; 2: UserDef {0-2}
  parameter PORT_USERDEF_ENABLED      = 1,           // The User-Defined port is visible to the customer {0,1}
  parameter PORT_ERR_RESP_ENABLED     = 0,           // The Errored Response port is visible to the customer {0,1}
  parameter TX_ENABLE_FAIRNESS        = 1)           // If set, I/O can be rerouted to the maint port {0,1}
  // }}} end LOG Parameters
(
  // {{{ Port Declarations -----------------
  // System Interface
  //----------------------------------------
  input             log_clk,                 // LOG interface clock
  input             log_rst,                 // Reset for LOG clock Domain
  input             cfg_clk,                 // CFG Interface user clock
  input             cfg_rst,                 // Reset for CFG clk domain
  input             maintr_rst,              // Reset for maintr interface, on LOG clk domain

  // PORT A Inteface
  //----------------------------------------
  // Request Interface
  input             UG_tx_porta_tvalid,      // Indicates Valid Input on the Request Channel
  output            LA_tx_porta_tready,      // Beat has been accepted
  input             UG_tx_porta_tlast,       // Indicates last beat
  input  [63:0]     UG_tx_porta_tdata,       // Req Data Bus
  input  [7:0]      UG_tx_porta_tkeep,       // Req Keep Bus
  input  [39:0]     UG_tx_porta_tuser,       // Req User Bus

  // Response Interface
  output            LA_rx_porta_tvalid,      // Indicates Valid Output on the Response Channel
  input             UG_rx_porta_tready,      // Beat has been accepted
  output            LA_rx_porta_tlast,       // Indicates last beat
  output  [63:0]    LA_rx_porta_tdata,       // Resp Data Bus
  output  [7:0]     LA_rx_porta_tkeep,       // Resp Keep Bus
  output  [39:0]    LA_rx_porta_tuser,       // Resp User Bus

  // PORT B Inteface
  //----------------------------------------
  // Request Interface
  input             UG_tx_portb_tvalid,      // Indicates Valid Input on the Request Channel
  output            LA_tx_portb_tready,      // Beat has been accepted
  input             UG_tx_portb_tlast,       // Indicates last beat
  input  [63:0]     UG_tx_portb_tdata,       // Req Data Bus
  input  [7:0]      UG_tx_portb_tkeep,       // Req keep Bus
  input  [39:0]     UG_tx_portb_tuser,       // Req User Bus

  // Response Interface
  output            LA_rx_portb_tvalid,      // Indicates Valid Output on the Response Channel
  input             UG_rx_portb_tready,      // Beat has been accepted
  output            LA_rx_portb_tlast,       // Indicates last beat
  output  [63:0]    LA_rx_portb_tdata,       // Resp Data Bus
  output  [7:0]     LA_rx_portb_tkeep,       // Resp Keep Bus
  output  [39:0]    LA_rx_portb_tuser,       // Resp User Bus

  // PORT C Inteface
  //----------------------------------------
  // Request Interface
  input             UG_tx_portc_tvalid,      // Indicates Valid Input on the Request Channel
  output            LA_tx_portc_tready,      // Beat has been accepted
  input             UG_tx_portc_tlast,       // Indicates last beat
  input  [63:0]     UG_tx_portc_tdata,       // Req Data Bus
  input  [7:0]      UG_tx_portc_tkeep,       // Req Keep Bus
  input  [39:0]     UG_tx_portc_tuser,       // Req User Bus

  // Response Interface
  output            LA_rx_portc_tvalid,      // Indicates Valid Output on the Response Channel
  input             UG_rx_portc_tready,      // Beat has been accepted
  output            LA_rx_portc_tlast,       // Indicates last beat
  output  [63:0]    LA_rx_portc_tdata,       // Resp Data Bus
  output  [7:0]     LA_rx_portc_tkeep,       // Resp Keep Bus
  output  [39:0]    LA_rx_portc_tuser,       // Resp User Bus

  // PORT D Inteface
  //----------------------------------------
  // Request Interface
  input             UG_tx_portd_tvalid,      // Indicates Valid Input on the Request Channel
  output            LA_tx_portd_tready,      // Beat has been accepted
  input             UG_tx_portd_tlast,       // Indicates last beat
  input  [63:0]     UG_tx_portd_tdata,       // Req Data Bus
  input  [7:0]      UG_tx_portd_tkeep,       // Req Keep Bus
  input  [39:0]     UG_tx_portd_tuser,       // Req User Bus

  // Response Interface
  output            LA_rx_portd_tvalid,      // Indicates Valid Output on the Response Channel
  input             UG_rx_portd_tready,      // Beat has been accepted
  output            LA_rx_portd_tlast,       // Indicates last beat
  output  [63:0]    LA_rx_portd_tdata,       // Resp Data Bus
  output  [7:0]     LA_rx_portd_tkeep,       // Resp Keep Bus
  output  [39:0]    LA_rx_portd_tuser,       // Resp User Bus

  // PORT E Inteface
  //----------------------------------------
  // Request Interface
  input             UG_tx_porte_tvalid,      // Indicates Valid Input on the Request Channel
  output            LA_tx_porte_tready,      // Beat has been accepted
  input             UG_tx_porte_tlast,       // Indicates last beat
  input  [63:0]     UG_tx_porte_tdata,       // Req Data Bus
  input  [7:0]      UG_tx_porte_tkeep,       // Req Keep Bus
  input  [39:0]     UG_tx_porte_tuser,       // Req User Bus

  // Response Interface
  output            LA_rx_porte_tvalid,      // Indicates Valid Output on the Response Channel
  input             UG_rx_porte_tready,      // Beat has been accepted
  output            LA_rx_porte_tlast,       // Indicates last beat
  output  [63:0]    LA_rx_porte_tdata,       // Resp Data Bus
  output  [7:0]     LA_rx_porte_tkeep,       // Resp Keep Bus
  output  [39:0]    LA_rx_porte_tuser,       // Resp User Bus

  // PORT F Inteface
  //----------------------------------------
  // Request Interface
  input             UG_tx_portf_tvalid,      // Indicates Valid Input on the Request Channel
  output            LA_tx_portf_tready,      // Beat has been accepted
  input             UG_tx_portf_tlast,       // Indicates last beat
  input  [63:0]     UG_tx_portf_tdata,       // Req Data Bus
  input  [7:0]      UG_tx_portf_tkeep,       // Req Keep Bus
  input  [39:0]     UG_tx_portf_tuser,       // Req User Bus

  // Response Interface
  output            LA_rx_portf_tvalid,      // Indicates Valid Output on the Response Channel
  input             UG_rx_portf_tready,      // Beat has been accepted
  output            LA_rx_portf_tlast,       // Indicates last beat
  output  [63:0]    LA_rx_portf_tdata,       // Resp Data Bus
  output  [7:0]     LA_rx_portf_tkeep,       // Resp Keep Bus
  output  [39:0]    LA_rx_portf_tuser,       // Resp User Bus

  // PORT G Inteface
  //----------------------------------------
  // Request Interface
  input             UG_tx_portg_tvalid,      // Indicates Valid Input on the Request Channel
  output            LA_tx_portg_tready,      // Beat has been accepted
  input             UG_tx_portg_tlast,       // Indicates last beat
  input  [63:0]     UG_tx_portg_tdata,       // Req Data Bus
  input  [7:0]      UG_tx_portg_tkeep,       // Req Keep Bus
  input  [39:0]     UG_tx_portg_tuser,       // Req User Bus

  // Response Interface
  output            LA_rx_portg_tvalid,      // Indicates Valid Output on the Response Channel
  input             UG_rx_portg_tready,      // Beat has been accepted
  output            LA_rx_portg_tlast,       // Indicates last beat
  output  [63:0]    LA_rx_portg_tdata,       // Resp Data Bus
  output  [7:0]     LA_rx_portg_tkeep,       // Resp keep Bus
  output  [39:0]    LA_rx_portg_tuser,       // Resp User Bus

  // PORT H Inteface
  //----------------------------------------
  // Request Interface
  input             UG_tx_porth_tvalid,      // Indicates Valid Input on the Request Channel
  output            LA_tx_porth_tready,      // Beat has been accepted
  input             UG_tx_porth_tlast,       // Indicates last beat
  input  [63:0]     UG_tx_porth_tdata,       // Req Data Bus
  input  [7:0]      UG_tx_porth_tkeep,       // Req Keep Bus
  input  [39:0]     UG_tx_porth_tuser,       // Req User Bus

  // Response Interface
  output            LA_rx_porth_tvalid,      // Indicates Valid Output on the Response Channel
  input             UG_rx_porth_tready,      // Beat has been accepted
  output            LA_rx_porth_tlast,       // Indicates last beat
  output  [63:0]    LA_rx_porth_tdata,       // Resp Data Bus
  output  [7:0]     LA_rx_porth_tkeep,       // Resp Keep Bus
  output  [39:0]    LA_rx_porth_tuser,       // Resp User Bus

  // Maintenance Interface
  //----------------------------------------
  input              UG_maintr_awvalid,      // Write Command Valid
  output             LR_maintr_awready,      // Write Port Ready
  input  [31:0]      UG_maintr_awaddr,       // Write Address
  input              UG_maintr_wvalid,       // Write Data Valid
  output             LR_maintr_wready,       // Write Port Ready
  input  [31:0]      UG_maintr_wdata,        // Write Data
  output             LR_maintr_bvalid,       // Write Response Valid
  input              UG_maintr_bready,       // Write Response Fabric Ready
  output [1:0]       LR_maintr_bresp,        // Write Response

  input              UG_maintr_arvalid,      // Read Command Valid
  output             LR_maintr_arready,      // Read Port Ready
  input  [31:0]      UG_maintr_araddr,       // Read Address
  output             LR_maintr_rvalid,       // Read Response Valid
  input              UG_maintr_rready,       // Read Response Fabric Ready
  output [31:0]      LR_maintr_rdata,        // Read Data
  output [1:0]       LR_maintr_rresp,        // Read Response


  // Maintenace/Config Fabric Interface
  //----------------------------------------
  // Write Request Port
  output            LR_cfgr_awvalid,         // Write Command Valid
  input             CF_cfgr_awready,         // Write Port Ready
  output [23:0]     LR_cfgr_awaddr,          // Write Address
  output            LR_cfgr_wvalid,          // Write Data Valid
  input             CF_cfgr_wready,          // Write Port Ready
  output [31:0]     LR_cfgr_wdata,           // Write Data
  output [3:0]      LR_cfgr_wstrb,           // Write Data byte enables
  output [2:0]      LR_cfgr_awprot,          // Write Protection (Tied to 0)

  // Write Response Port
  input             CF_cfgr_bvalid,          // Write Response Valid
  output            LR_cfgr_bready,          // Write Response Fabric Ready
  input  [1:0]      CF_cfgr_bresp,           // Write Response

  // Read Request Port
  output            LR_cfgr_arvalid,         // Read Command Valid
  input             CF_cfgr_arready,         // Read Port Ready
  output [23:0]     LR_cfgr_araddr,          // Read Address
  output [2:0]      LR_cfgr_arprot,          // Read Protection (Tied to 0)

  // Read Resposne Port
  input             CF_cfgr_rvalid,          // Read Response Valid
  output            LR_cfgr_rready,          // Read Response Fabric Ready
  input  [31:0]     CF_cfgr_rdata,           // Read Data
  input  [1:0]      CF_cfgr_rresp,           // Read Response

  // LOG/Buffer TX Interface
  //----------------------------------------
  output            LD_buft_tvalid,          // Valid packet beat
  input             BT_buft_tready,          // Packet beat accepted
  output [63:0]     LD_buft_tdata,           // Packet data
  output [7:0]      LD_buft_tkeep,           // Valid bytes in this beat, only valid on last
  output            LD_buft_tlast,           // Last beat
  output [7:0]      LD_buft_tuser,           // {4'h00, Response, VC, CRF, 1'b0}

  // Sideband
  input             BT_response_only,        // Disable requests

  // LOG/Buffer RX Interface
  //----------------------------------------
  input             BR_bufr_tvalid,          // Valid packet beat
  output            LE_bufr_tready,          // Packet beat accepted
  input  [63:0]     BR_bufr_tdata,           // Packet data
  input  [7:0]      BR_bufr_tkeep,           // Valid bytes in this beat, only valid on last
  input             BR_bufr_tlast,           // Last beat
  input  [7:0]      BR_bufr_tuser,           // {5'h00, VC, CRF, 1'b0}

  // Config Fabric to LOG CFG Registers Interface
  //----------------------------------------
  input             CF_cfgl_awvalid,         // Write Command Valid
  output            LC_cfgl_awready,         // Write Port Ready
  input  [23:0]     CF_cfgl_awaddr,          // Write Address
  input             CF_cfgl_wvalid,          // Write Data Valid
  output            LC_cfgl_wready,          // Write Port Ready
  input  [31:0]     CF_cfgl_wdata,           // Write Data
  input  [3:0]      CF_cfgl_wstrb,           // Write Data byte enables
  output            LC_cfgl_bvalid,          // Write Response Valid
  input             CF_cfgl_bready,          // Write Response Fabric Ready
  input             CF_cfgl_arvalid,         // Read Command Valid
  output            LC_cfgl_arready,         // Read Port Ready
  input  [23:0]     CF_cfgl_araddr,          // Read Address
  output            LC_cfgl_rvalid,          // Read Response Valid
  input             CF_cfgl_rready,          // Read Response Fabric Ready
  output [31:0]     LC_cfgl_rdata,           // Read Data

  //Sideband
  output [15:0]     LC_deviceid,             // Current DeviceID from the DeviceID register
  input             PC_maint_only,           // LOG can only send maint transactions
  output            LA_port_decode_error     // No valid output port for the RX transaction
  // }}} end port declarations -------------
);

// added below macro to fix the CR# 735137
// synthesis translate_off 
  // {{{ Invalid Parameter Checks
  initial begin
    if (PORT_ERR_RESP_ENABLED && (PORT_IO_STYLE != 2)) begin
      $display("ERROR: The error port cannot be enabled with PORT_IO_STYLE==%0d",PORT_IO_STYLE);
      $finish;
    end
    if (PORT_MAINT_STYLE == 0) begin
      $display("ERROR: Maintenance transaction can not be configured to use the IO ports.");
      $finish;
    end
    if (PORT_MAINT_STYLE == 2 && PORT_USERDEF_ENABLED == 0) begin
      $display("ERROR: Maintenance transactions were configured to use the USERDEF port, but the USERDEF port was not enabled.");
      $finish;
    end
  end
  // }}} end Invalid Parameter Checks
// synthesis translate_on

  //  {{{ Parameter Configuration
  //  + {{{ Arb TX Parameter Configuration +
  // Specify whether each port uses HELLO format {0,1}
  localparam TX_PORTA_HELLO             = PORT_IO_HELLO && !PORT_USERDEF_ENABLED;
  localparam TX_PORTB_HELLO             = PORT_IO_HELLO;
  localparam TX_PORTC_HELLO             = PORT_IO_HELLO;
  localparam TX_PORTD_HELLO             = PORT_IO_HELLO;
  localparam TX_PORTE_HELLO             = PORT_MSG_HELLO;
  localparam TX_PORTF_HELLO             = PORT_MSG_HELLO;
  localparam TX_PORTG_HELLO             = PORT_MAINT_HELLO;
  localparam TX_PORTH_HELLO             = PORT_MAINT_HELLO;

  // Specify whether each port is enabled
  localparam TX_PORTA_ENABLE            = (PORT_IO_STYLE > 1) || PORT_USERDEF_ENABLED;
  localparam TX_PORTB_ENABLE            = (PORT_IO_STYLE > 1);
  localparam TX_PORTC_ENABLE            = (PORT_IO_STYLE > 0);
  localparam TX_PORTD_ENABLE            = 1;
  localparam TX_PORTE_ENABLE            = (PORT_MSG_STYLE   == 1);
  localparam TX_PORTF_ENABLE            = (PORT_MSG_STYLE   == 1);
  localparam TX_PORTG_ENABLE            = (PORT_MAINT_STYLE == 1);
  localparam TX_PORTH_ENABLE            = (PORT_MAINT_STYLE == 1);

  // Per-port arbitration priority {0, 1, 2, 3}
  localparam TX_PORTA_PRIORITY          = 1;
  localparam TX_PORTB_PRIORITY          = 1;
  localparam TX_PORTC_PRIORITY          = 1;
  localparam TX_PORTD_PRIORITY          = 1;
  localparam TX_PORTE_PRIORITY          = 1;
  localparam TX_PORTF_PRIORITY          = 1;
  localparam TX_PORTG_PRIORITY          = 1;
  localparam TX_PORTH_PRIORITY          = 1;

  // Specify whether port is dedicated to response packets
  localparam TX_PORTA_RESP_CLASS        = 0; // User-Def TX or Read Initiator Request Port
  localparam TX_PORTB_RESP_CLASS        = 1; // Read Target Response Port
  localparam TX_PORTC_RESP_CLASS        = 0; // Initiator Request or Write Initiator Request Port
  localparam TX_PORTD_RESP_CLASS        = 1; // I/O or Target Response or Write Target Response Port
  localparam TX_PORTE_RESP_CLASS        = 0; // Msg Request Port
  localparam TX_PORTF_RESP_CLASS        = 1; // Msg Response Port
  localparam TX_PORTG_RESP_CLASS        = 0; // Maint Request Port
  localparam TX_PORTH_RESP_CLASS        = 1; // Maint Response Port
  //  + }}} end Arb TX Parameter Configuration +

  //  + {{{ Arb RX Parameter Configuration +
  // RX_PORTx_ENABLE_FTYPE_SORT  - 7-bit mask of FTYPEs to search for
  // RX_PORTx_FTYPE_SORT1        - FTYPE search pattern 1
  // RX_PORTx_FTYPE_SORT2        - FTYPE search pattern 2
  // RX_PORTx_FTYPE_SORT3        - FTYPE search pattern 3
  // RX_PORTx_FTYPE_SORT4        - FTYPE search pattern 4
  // RX_PORTx_FTYPE_SORT5        - FTYPE search pattern 5
  // RX_PORTx_FTYPE_SORT6        - FTYPE search pattern 6
  // RX_PORTx_FTYPE_SORT7        - FTYPE search pattern 7
  // RX_PORTx_ENABLE_TTYPE_SORT  - 7-bit mask of TTYPEs to search for (must also have corresponding FTYPE_SORT set)
  // RX_PORTx_TTYPE_SORT1        - TTYPE search pattern 1
  // RX_PORTx_TTYPE_SORT2        - TTYPE search pattern 2
  // RX_PORTx_TTYPE_SORT3        - TTYPE search pattern 3
  // RX_PORTx_TTYPE_SORT4        - TTYPE search pattern 4
  // RX_PORTx_TTYPE_SORT5        - TTYPE search pattern 5
  // RX_PORTx_TTYPE_SORT6        - TTYPE search pattern 6
  // RX_PORTx_TTYPE_SORT7        - TTYPE search pattern 7
  // RX_PORTx_ENABLE_STAT_SORT   - how many different STATs to look for {0-2}
  // RX_PORTx_STAT_SORT1         - STAT search pattern 1
  // RX_PORTx_STAT_SORT2         - STAT search pattern 2
  // RX_PORTx_LCSBA_SUPPORT      - If set, pkts will be routed to this port if the address matches the LCSBA mask {0,1}

  localparam INIT_MSG                   = ((MSG_INIT_SINGLE == 1) || (MSG_INIT_MULTI == 1));
  localparam TARGET_MSG                 = ((MSG_SINK_SINGLE == 1) || (MSG_SINK_MULTI == 1));

  localparam [3:0] FTYPE_NREAD          = 4'b0010;
  localparam [3:0] FTYPE_NWRITE         = 4'b0101;
  localparam [3:0] FTYPE_SWRITE         = 4'b0110;
  localparam [3:0] FTYPE_MAINT          = 4'b1000;
  localparam [3:0] FTYPE_DS             = 4'b1001;
  localparam [3:0] FTYPE_DB             = 4'b1010;
  localparam [3:0] FTYPE_MSG            = 4'b1011;
  localparam [3:0] FTYPE_RESP           = 4'b1101;
  localparam [3:0] TTYPE_MAINT_RREQ     = 4'b0000;
  localparam [3:0] TTYPE_MAINT_WREQ     = 4'b0001;
  localparam [3:0] TTYPE_MAINT_RRESP    = 4'b0010;
  localparam [3:0] TTYPE_MAINT_WRESP    = 4'b0011;
  localparam [3:0] TTYPE_RESP_NODATA    = 4'b0000;
  localparam [3:0] TTYPE_RESP_WDATA     = 4'b1000;
  localparam [3:0] TTYPE_RESP_MSG       = 4'b0001;
  localparam [3:0] RESP_STATUS_ERR      = 4'b0111;
  localparam [3:0] RESP_STATUS_DONE     = 4'b0000;

  // RX Port A Configuration
  // -----------------------
  // RX Port A is the Read Initiator Response port if in Independent Read/Write
  // mode, otherwise it is the user-defined port (if enabled)
                                          // If set, unmatched pkts fall through to Porta {0,1}
  localparam RX_PORTA_FALL_THROUGH      = (PORT_IO_STYLE < 2) && PORT_USERDEF_ENABLED;
  localparam RX_PORTA_ENABLE_FTYPE_SORT =
               {6'b0, ((PORT_IO_STYLE == 2) && ((INIT_NREAD == 1) || (INIT_ATOMIC == 1)))};
  localparam RX_PORTA_FTYPE_SORT1       = FTYPE_RESP;
  localparam RX_PORTA_FTYPE_SORT2       = FTYPE_MAINT;
  localparam RX_PORTA_FTYPE_SORT3       = FTYPE_MAINT;
  localparam RX_PORTA_FTYPE_SORT4       = 1;
  localparam RX_PORTA_FTYPE_SORT5       = 1;
  localparam RX_PORTA_FTYPE_SORT6       = 1;
  localparam RX_PORTA_FTYPE_SORT7       = 1;
  localparam RX_PORTA_ENABLE_TTYPE_SORT =
               {6'b0, ((PORT_IO_STYLE == 2) && ((INIT_NREAD == 1) || (INIT_ATOMIC == 1)))};
  localparam RX_PORTA_TTYPE_SORT1       = TTYPE_RESP_WDATA;
  localparam RX_PORTA_TTYPE_SORT2       = 1;
  localparam RX_PORTA_TTYPE_SORT3       = 1;
  localparam RX_PORTA_TTYPE_SORT4       = 1;
  localparam RX_PORTA_TTYPE_SORT5       = 1;
  localparam RX_PORTA_TTYPE_SORT6       = 1;
  localparam RX_PORTA_TTYPE_SORT7       = 1;
  localparam RX_PORTA_ENABLE_STAT_SORT  = 0;
  localparam RX_PORTA_STAT_SORT1        = 1;
  localparam RX_PORTA_STAT_SORT2        = 1;
  localparam RX_PORTA_LCSBA_SUPPORT     = 0;

  // RX Port B Configuration
  // -----------------------
  // RX Port B is the Read Target Request port if in Independent Read/Write
  // mode, otherwise it is unused
  localparam RX_PORTB_ENABLE_FTYPE_SORT = {5'b0, (PORT_MAINT_STYLE == 0), (PORT_IO_STYLE == 2)};
  localparam RX_PORTB_FTYPE_SORT1       = FTYPE_NREAD;
  localparam RX_PORTB_FTYPE_SORT2       = FTYPE_MAINT;
  localparam RX_PORTB_FTYPE_SORT3       = 1;
  localparam RX_PORTB_FTYPE_SORT4       = 1;
  localparam RX_PORTB_FTYPE_SORT5       = 1;
  localparam RX_PORTB_FTYPE_SORT6       = 1;
  localparam RX_PORTB_FTYPE_SORT7       = 1;
  localparam RX_PORTB_ENABLE_TTYPE_SORT = {5'b0, (PORT_MAINT_STYLE == 0), 1'b0};
  localparam RX_PORTB_TTYPE_SORT1       = 1;
  localparam RX_PORTB_TTYPE_SORT2       = TTYPE_MAINT_RREQ;
  localparam RX_PORTB_TTYPE_SORT3       = 1;
  localparam RX_PORTB_TTYPE_SORT4       = 1;
  localparam RX_PORTB_TTYPE_SORT5       = 1;
  localparam RX_PORTB_TTYPE_SORT6       = 1;
  localparam RX_PORTB_TTYPE_SORT7       = 1;
  localparam RX_PORTB_ENABLE_STAT_SORT  = 0;
  localparam RX_PORTB_STAT_SORT1        = 1;
  localparam RX_PORTB_STAT_SORT2        = 1;
  localparam RX_PORTB_LCSBA_SUPPORT     = 0;

  // RX Port C Configuration
  // -----------------------
  // RX Port C is the Initiator Response Port or the Write Initiator Response
  // Port, depending on I/O style.
  localparam RX_PORTC_ENABLE_FTYPE_SORT =
             {4'b0,
              // Messaging
              (((MSG_INIT_SINGLE == 1) || (MSG_INIT_MULTI == 1)) && (PORT_MSG_STYLE == 0) && (PORT_IO_STYLE > 0)),
              // Read Responses
              ((INIT_NREAD == 1) || (INIT_ATOMIC == 1)) && (PORT_IO_STYLE == 1),
              // Write Responses
              ((INIT_NWRITE_R == 1) || (INIT_DB == 1)) && (PORT_IO_STYLE > 0)};

  localparam RX_PORTC_FTYPE_SORT1       = FTYPE_RESP;
  localparam RX_PORTC_FTYPE_SORT2       = FTYPE_RESP;
  localparam RX_PORTC_FTYPE_SORT3       = FTYPE_RESP;
  localparam RX_PORTC_FTYPE_SORT4       = 1;
  localparam RX_PORTC_FTYPE_SORT5       = 1;
  localparam RX_PORTC_FTYPE_SORT6       = 1;
  localparam RX_PORTC_FTYPE_SORT7       = 1;

  localparam RX_PORTC_ENABLE_TTYPE_SORT =
             {4'b0,
              // Messaging
              (((MSG_INIT_SINGLE == 1) || (MSG_INIT_MULTI == 1)) && (PORT_MSG_STYLE == 0) && (PORT_IO_STYLE > 0)),
              // Read Responses
              ((INIT_NREAD == 1) || (INIT_ATOMIC == 1)) && (PORT_IO_STYLE == 1),
              // Write Responses
              ((INIT_NWRITE_R == 1) || (INIT_DB == 1)) && (PORT_IO_STYLE > 0)};

  localparam RX_PORTC_TTYPE_SORT1       = TTYPE_RESP_NODATA;
  localparam RX_PORTC_TTYPE_SORT2       = TTYPE_RESP_WDATA;
  localparam RX_PORTC_TTYPE_SORT3       = TTYPE_RESP_MSG;
  localparam RX_PORTC_TTYPE_SORT4       = 1;
  localparam RX_PORTC_TTYPE_SORT5       = 1;
  localparam RX_PORTC_TTYPE_SORT6       = 1;
  localparam RX_PORTC_TTYPE_SORT7       = 1;
  localparam RX_PORTC_ENABLE_STAT_SORT  = 0;
  localparam RX_PORTC_STAT_SORT1        = 1;
  localparam RX_PORTC_STAT_SORT2        = 1;
  localparam RX_PORTC_LCSBA_SUPPORT     = 0;

  // RX Port D Configuration
  // -----------------------
  // RX Port D is the Generic I/O port or the Target Request Port or the Write
  // Target Request Port, depending on I/O style.
  localparam RX_PORTD_ENABLE_FTYPE_SORT = {((PORT_MSG_STYLE < 1) && (TARGET_MSG      == 1)),
                                            (PORT_IO_STYLE <  1),
                                            (PORT_IO_STYLE <  1),
                                            (TARGET_DB     == 1),
                                            (TARGET_SWRITE == 1),
                                           ((TARGET_NWRITE == 1) || (TARGET_NWRITE_R == 1) || (TARGET_ATOMIC == 1)),
                                           ((PORT_IO_STYLE <  2) && ((TARGET_NREAD   == 1) || (TARGET_ATOMIC == 1)))};
  localparam RX_PORTD_FTYPE_SORT1       = FTYPE_NREAD;
  localparam RX_PORTD_FTYPE_SORT2       = FTYPE_NWRITE;
  localparam RX_PORTD_FTYPE_SORT3       = FTYPE_SWRITE;
  localparam RX_PORTD_FTYPE_SORT4       = FTYPE_DB;
  localparam RX_PORTD_FTYPE_SORT5       = FTYPE_RESP;
  localparam RX_PORTD_FTYPE_SORT6       = FTYPE_RESP;
  localparam RX_PORTD_FTYPE_SORT7       = FTYPE_MSG;
  localparam RX_PORTD_ENABLE_TTYPE_SORT = {1'b0, (PORT_MSG_STYLE > 0), (PORT_MSG_STYLE > 0), 4'b0};
  localparam RX_PORTD_TTYPE_SORT1       = 1;
  localparam RX_PORTD_TTYPE_SORT2       = 1;
  localparam RX_PORTD_TTYPE_SORT3       = 1;
  localparam RX_PORTD_TTYPE_SORT4       = 1;
  localparam RX_PORTD_TTYPE_SORT5       = TTYPE_RESP_NODATA;
  localparam RX_PORTD_TTYPE_SORT6       = TTYPE_RESP_WDATA;
  localparam RX_PORTD_TTYPE_SORT7       = 1;
  localparam RX_PORTD_ENABLE_STAT_SORT  = 0;
  localparam RX_PORTD_STAT_SORT1        = 1;
  localparam RX_PORTD_STAT_SORT2        = 1;
  localparam RX_PORTD_LCSBA_SUPPORT     = 0;

  // RX Port E Configuration
  // -----------------------
  // RX Port E is the Message Initiator Response port if it exists.
  localparam RX_PORTE_ENABLE_FTYPE_SORT = {6'b0, (PORT_MSG_STYLE == 1)};
  localparam RX_PORTE_FTYPE_SORT1       = FTYPE_RESP;
  localparam RX_PORTE_FTYPE_SORT2       = 1;
  localparam RX_PORTE_FTYPE_SORT3       = 1;
  localparam RX_PORTE_FTYPE_SORT4       = 1;
  localparam RX_PORTE_FTYPE_SORT5       = 1;
  localparam RX_PORTE_FTYPE_SORT6       = 1;
  localparam RX_PORTE_FTYPE_SORT7       = 1;
  localparam RX_PORTE_ENABLE_TTYPE_SORT = {6'b0, (PORT_MSG_STYLE == 1)};
  localparam RX_PORTE_TTYPE_SORT1       = TTYPE_RESP_MSG;
  localparam RX_PORTE_TTYPE_SORT2       = 1;
  localparam RX_PORTE_TTYPE_SORT3       = 1;
  localparam RX_PORTE_TTYPE_SORT4       = 1;
  localparam RX_PORTE_TTYPE_SORT5       = 1;
  localparam RX_PORTE_TTYPE_SORT6       = 1;
  localparam RX_PORTE_TTYPE_SORT7       = 1;
  localparam RX_PORTE_ENABLE_STAT_SORT  = 0;
  localparam RX_PORTE_STAT_SORT1        = 1;
  localparam RX_PORTE_STAT_SORT2        = 1;
  localparam RX_PORTE_LCSBA_SUPPORT     = 0;

  // RX Port F Configuration
  // -----------------------
  // RX Port F is the Message Target Request port if it exists.
  localparam RX_PORTF_ENABLE_FTYPE_SORT = {6'b0,(PORT_MSG_STYLE == 1)};
  localparam RX_PORTF_FTYPE_SORT1       = FTYPE_MSG;
  localparam RX_PORTF_FTYPE_SORT2       = 1;
  localparam RX_PORTF_FTYPE_SORT3       = 1;
  localparam RX_PORTF_FTYPE_SORT4       = 1;
  localparam RX_PORTF_FTYPE_SORT5       = 1;
  localparam RX_PORTF_FTYPE_SORT6       = 1;
  localparam RX_PORTF_FTYPE_SORT7       = 1;
  localparam RX_PORTF_ENABLE_TTYPE_SORT = 0;
  localparam RX_PORTF_TTYPE_SORT1       = 1;
  localparam RX_PORTF_TTYPE_SORT2       = 1;
  localparam RX_PORTF_TTYPE_SORT3       = 1;
  localparam RX_PORTF_TTYPE_SORT4       = 1;
  localparam RX_PORTF_TTYPE_SORT5       = 1;
  localparam RX_PORTF_TTYPE_SORT6       = 1;
  localparam RX_PORTF_TTYPE_SORT7       = 1;
  localparam RX_PORTF_ENABLE_STAT_SORT  = 0;
  localparam RX_PORTF_STAT_SORT1        = 1;
  localparam RX_PORTF_STAT_SORT2        = 1;
  localparam RX_PORTF_LCSBA_SUPPORT     = 0;

  // RX Port G Configuration
  // -----------------------
  // RX Port G is the Errored Response port if it exists. Errored I/O responses
  // go here (both TTYPEs of response with data or response w/o data). If MSGs
  // are assigned to the I/O port, (PORT_MSG_STYLE=0), errored MSG responses go
  // here too.
  localparam RX_PORTG_ENABLE_FTYPE_SORT = {5'b0, {2{(PORT_ERR_RESP_ENABLED == 1)}} };
  localparam RX_PORTG_FTYPE_SORT1       = FTYPE_RESP;
  localparam RX_PORTG_FTYPE_SORT2       = FTYPE_RESP;
  localparam RX_PORTG_FTYPE_SORT3       = 1;
  localparam RX_PORTG_FTYPE_SORT4       = 1;
  localparam RX_PORTG_FTYPE_SORT5       = 1;
  localparam RX_PORTG_FTYPE_SORT6       = 1;
  localparam RX_PORTG_FTYPE_SORT7       = 1;
  localparam RX_PORTG_ENABLE_TTYPE_SORT = {5'b0, {2{(PORT_ERR_RESP_ENABLED == 1)}} };
  localparam RX_PORTG_TTYPE_SORT1       = TTYPE_RESP_NODATA;
  localparam RX_PORTG_TTYPE_SORT2       = TTYPE_RESP_WDATA;
  localparam RX_PORTG_TTYPE_SORT3       = 1;
  localparam RX_PORTG_TTYPE_SORT4       = 1;
  localparam RX_PORTG_TTYPE_SORT5       = 1;
  localparam RX_PORTG_TTYPE_SORT6       = 1;
  localparam RX_PORTG_TTYPE_SORT7       = 1;
  localparam RX_PORTG_ENABLE_STAT_SORT  = {1'b0, (PORT_ERR_RESP_ENABLED == 1)};
  localparam RX_PORTG_STAT_SORT1        = RESP_STATUS_ERR;
  localparam RX_PORTG_STAT_SORT2        = 1;
  localparam RX_PORTG_LCSBA_SUPPORT     = 0;

  // RX Port H Configuration
  // -----------------------
  // RX Port H is the Maintenance port if it exists. All MAINT transactions go
  // here (requests and responses).
  localparam RX_PORTH_ENABLE_FTYPE_SORT = {6'b0, (PORT_MAINT_STYLE == 1)};
  localparam RX_PORTH_FTYPE_SORT1       = FTYPE_MAINT;
  localparam RX_PORTH_FTYPE_SORT2       = 1;
  localparam RX_PORTH_FTYPE_SORT3       = 1;
  localparam RX_PORTH_FTYPE_SORT4       = 1;
  localparam RX_PORTH_FTYPE_SORT5       = 1;
  localparam RX_PORTH_FTYPE_SORT6       = 1;
  localparam RX_PORTH_FTYPE_SORT7       = 1;
  localparam RX_PORTH_ENABLE_TTYPE_SORT = 0;
  localparam RX_PORTH_TTYPE_SORT1       = 1;
  localparam RX_PORTH_TTYPE_SORT2       = 1;
  localparam RX_PORTH_TTYPE_SORT3       = 1;
  localparam RX_PORTH_TTYPE_SORT4       = 1;
  localparam RX_PORTH_TTYPE_SORT5       = 1;
  localparam RX_PORTH_TTYPE_SORT6       = 1;
  localparam RX_PORTH_TTYPE_SORT7       = 1;
  localparam RX_PORTH_ENABLE_STAT_SORT  = 0;
  localparam RX_PORTH_STAT_SORT1        = 1;
  localparam RX_PORTH_STAT_SORT2        = 1;
  localparam RX_PORTH_LCSBA_SUPPORT     = LCSBA_SUPPORT;
  //  + }}} end Arb RX Parameter Configuration +

  //  + {{{ HELLO Decoder Parameter Configuration +
  localparam DECODE_FT02                = (PORT_IO_HELLO    == 1) && ((INIT_NREAD   == 1)    || (INIT_ATOMIC == 1));
  localparam DECODE_FT05                = (PORT_IO_HELLO    == 1) &&
                                         ((INIT_NWRITE      == 1) ||  (INIT_NWRITE_R == 1)   || (INIT_ATOMIC == 1));
  localparam DECODE_FT06                = (PORT_IO_HELLO    == 1) &&  (INIT_SWRITE   == 1);
  localparam DECODE_FT08                = (PORT_MAINT_HELLO == 1) &&  (MAINT_SOURCE  == 1);
  localparam DECODE_FT09                = (PORT_IO_HELLO    == 1) &&  (INIT_DS       == 1);
  localparam DECODE_FT10                = (PORT_IO_HELLO    == 1) &&  (INIT_DB       == 1);
  localparam DECODE_FT11                = (PORT_MSG_HELLO   == 1) && ((MSG_INIT_SINGLE == 1) || (MSG_INIT_MULTI == 1));
  localparam DECODE_FT13                = (PORT_IO_HELLO    == 1) ||  (PORT_MSG_HELLO   == 1);
  //  + }}} HELLO Decoder Parameter Configuration +
  //  }}} end Parameter Configuration

  // {{{ Between the Arb and CFG
  wire [9:0]            LC_lcsba;               // Local Configuration Space Base Address msbs
  // }}}

  // {{{ Between the Maint and Arb
  // TX Request Interface
  //----------------------------------------
  wire                  LR_lrtx_req_tvalid;     // Valid packet beat
  wire                  LA_lrtx_req_tready;     // Packet beat accepted
  wire       [63:0]     LR_lrtx_req_tdata;      // Packet data
  wire       [7:0]      LR_lrtx_req_tkeep;      // Valid bytes in this beat, only valid on last
  wire                  LR_lrtx_req_tlast;      // Last beat
  wire       [39:0]     LR_lrtx_req_tuser;      // {SrcID, DestID, 3'b0, Response (1'b0), 1'b0, CRF, 1'b0}

  // TX Response Interface
  //----------------------------------------
  wire                  LR_lrtx_resp_tvalid;    // Valid packet beat
  wire                  LA_lrtx_resp_tready;    // Packet beat accepted
  wire       [63:0]     LR_lrtx_resp_tdata;     // Packet data
  wire       [7:0]      LR_lrtx_resp_tkeep;     // Valid bytes in this beat, only valid on last
  wire                  LR_lrtx_resp_tlast;     // Last beat
  wire       [39:0]     LR_lrtx_resp_tuser;     // {SrcID, DestID, 3'b0, Response (1'b1), 1'b0, CRF, 1'b0}

  // RX Interface
  //----------------------------------------
  wire                  LA_lrrx_tvalid;         // Valid packet beat
  wire                  LR_lrrx_tready;         // Packet beat accepted
  wire       [63:0]     LA_lrrx_tdata;          // Packet data
  wire       [7:0]      LA_lrrx_tkeep;          // Valid bytes in this beat, only valid on last
  wire                  LA_lrrx_tlast;          // Last beat
  wire       [39:0]     LA_lrrx_tuser;          // {SrcID, DestID, 3'b0, Response, 1'b0, CRF, 1'b0}

  // TX Request Interface
  //----------------------------------------
  wire                  UG_tx_portg_tvalid_int; // Valid packet beat
  wire                  LA_tx_portg_tready_int; // Packet beat accepted
  wire       [63:0]     UG_tx_portg_tdata_int;  // Packet data
  wire       [7:0]      UG_tx_portg_tkeep_int;  // Valid bytes in this beat, only valid on last
  wire                  UG_tx_portg_tlast_int;  // Last beat
  wire       [39:0]     UG_tx_portg_tuser_int;  // {SrcID, DestID, 3'b0, Response (1'b0), 1'b0, CRF, 1'b0}

  // TX Response Interface
  //----------------------------------------
  wire                  UG_tx_porth_tvalid_int; // Valid packet beat
  wire                  LA_tx_porth_tready_int; // Packet beat accepted
  wire       [63:0]     UG_tx_porth_tdata_int;  // Packet data
  wire       [7:0]      UG_tx_porth_tkeep_int;  // Valid bytes in this beat, only valid on last
  wire                  UG_tx_porth_tlast_int;  // Last beat
  wire       [39:0]     UG_tx_porth_tuser_int;  // {SrcID, DestID, 3'b0, Response (1'b1), 1'b0, CRF, 1'b0}

  // RX Interface
  //----------------------------------------
  wire                  LA_rx_porth_tvalid_int; // Valid packet beat
  wire                  UG_rx_porth_tready_int; // Packet beat accepted
  wire       [63:0]     LA_rx_porth_tdata_int;  // Packet data
  wire       [7:0]      LA_rx_porth_tkeep_int;  // Valid bytes in this beat, only valid on last
  wire                  LA_rx_porth_tlast_int;  // Last beat
  wire       [39:0]     LA_rx_porth_tuser_int;  // {SrcID, DestID, 3'b0, Response, 1'b0, CRF, 1'b0}
  // }}}

  // {{{ Between the Arb and Encoder
  // RX Interface
  //----------------------------------------
  wire                  LE_lhrx_tvalid;         // Valid Packet Beat
  wire                  LA_lhrx_tready;         // Packet Beat Accepted
  wire       [63:0]     LE_lhrx_tdata;          // Packet Data
  wire        [7:0]     LE_lhrx_tkeep;          // Valid bytes in this beat, only valid on last
  wire                  LE_lhrx_tlast;          // Last Beat
  wire       [39:0]     LE_lhrx_tuser;          // {DEST_ID, SRC_ID, 2'h0, HELLO_FMT, 2'h0, VC, CRF, 1'b0}
  wire                  LE_unsupported_type;    // The packet has been decoded as an unsupported type

  // TX Interface
  //----------------------------------------
  wire                  LA_lhtx_tvalid;         // Valid Packet Beat
  wire                  LD_lhtx_tready;         // Packet Beat Accepted
  wire       [63:0]     LA_lhtx_tdata;          // Packet Data
  wire        [7:0]     LA_lhtx_tkeep;          // Valid bytes in this beat, only valid on last
  wire                  LA_lhtx_tlast;          // Last Beat
  wire       [39:0]     LA_lhtx_tuser;          // {DEST_ID, SRC_ID, 3'h0, RESPONSE, HELLO_FMT, VC, CRF, 1'b0}
  // }}}



  // {{{ log_cfg_top instantiation
  //----------------------------------------
  srio_gen2_v4_1_16_log_cfg_top
    #(.TCQ                       (TCQ),
      .HW_ARCH                   (HW_ARCH),
      .DEVICEID_WIDTH            (DEVICEID_WIDTH),
      .DEVICEID                  (DEVICEID),
      .INIT_NREAD                (INIT_NREAD),
      .INIT_NWRITE               (INIT_NWRITE),
      .INIT_SWRITE               (INIT_SWRITE),
      .INIT_NWRITE_R             (INIT_NWRITE_R),
      .INIT_DB                   (INIT_DB),
      .INIT_DS                   (INIT_DS),
      .INIT_ATOMIC               (INIT_ATOMIC),
      .MSG_INIT_SINGLE           (MSG_INIT_SINGLE),
      .MSG_INIT_MULTI            (MSG_INIT_MULTI),
      .TARGET_NREAD              (TARGET_NREAD),
      .TARGET_NWRITE             (TARGET_NWRITE),
      .TARGET_SWRITE             (TARGET_SWRITE),
      .TARGET_NWRITE_R           (TARGET_NWRITE_R),
      .TARGET_DB                 (TARGET_DB),
      .TARGET_DS                 (TARGET_DS),
      .TARGET_ATOMIC             (TARGET_ATOMIC),
      .MSG_SINK_SINGLE           (MSG_SINK_SINGLE),
      .MSG_SINK_MULTI            (MSG_SINK_MULTI),
      .CRF_SUPPORT               (CRF_SUPPORT),
      .DEVID_CAR                 (DEVID_CAR),
      .DEVINFO_CAR               (DEVINFO_CAR),
      .DEV_CAR_OVRD              (DEV_CAR_OVRD),
      .LCSBA_SUPPORT             (LCSBA_SUPPORT),
      .LCSBA                     (LCSBA),
      .ASSY_ID                   (ASSY_ID),
      .ASSY_VENDOR               (ASSY_VENDOR),
      .ASSY_REV                  (ASSY_REV),
      .PE_BRIDGE                 (PE_BRIDGE),
      .PE_MEMORY                 (PE_MEMORY),
      .PE_PROC                   (PE_PROC),
      .PE_SWITCH                 (PE_SWITCH),
      .PHY_EF_PTR                (PHY_EF_PTR))
    log_cfg_top_inst
     (.log_clk                   (log_clk),
      .log_rst                   (log_rst),
      .cfg_clk                   (cfg_clk),
      .cfg_rst                   (cfg_rst),
      .LC_deviceid               (LC_deviceid),
      .LC_lcsba                  (LC_lcsba),
      .CF_cfgl_awvalid           (CF_cfgl_awvalid),
      .LC_cfgl_awready           (LC_cfgl_awready),
      .CF_cfgl_awaddr            (CF_cfgl_awaddr),
      .CF_cfgl_wvalid            (CF_cfgl_wvalid),
      .LC_cfgl_wready            (LC_cfgl_wready),
      .CF_cfgl_wdata             (CF_cfgl_wdata),
      .CF_cfgl_wstrb             (CF_cfgl_wstrb),
      .LC_cfgl_bvalid            (LC_cfgl_bvalid),
      .CF_cfgl_bready            (CF_cfgl_bready),
      .CF_cfgl_arvalid           (CF_cfgl_arvalid),
      .LC_cfgl_arready           (LC_cfgl_arready),
      .CF_cfgl_araddr            (CF_cfgl_araddr),
      .LC_cfgl_rvalid            (LC_cfgl_rvalid),
      .CF_cfgl_rready            (CF_cfgl_rready),
      .LC_cfgl_rdata             (LC_cfgl_rdata)
     );
  // }}} End log_cfg_top instantiation

// Generate used to instantiate log_maint or not, depending on MAINT_CFG
// Aliasing of the signals is needed for the arbiter ports that the maint
// uses because ports can't be generated.
generate if (MAINT_CFG == 1) begin: maint_block_enabled_gen
  // {{{ log_maint instantiation
  //--------------------------------------------
  srio_gen2_v4_1_16_log_maint
    #(.TCQ                       (TCQ),
      .DEVICEID_WIDTH            (DEVICEID_WIDTH),
      .TARGET_NREAD              (TARGET_NREAD),
      .TARGET_NWRITE             (TARGET_NWRITE),
      .TARGET_NWRITE_R           (TARGET_NWRITE_R),
      .CRF_SUPPORT               (CRF_SUPPORT),
      .MAINT_SOURCE              (MAINT_SOURCE),
      .LCSBA_SUPPORT             (LCSBA_SUPPORT),
      .VC                        (VC))
    log_maint_inst
     (.log_clk                   (log_clk),
      .log_rst                   (log_rst),
      .maintr_rst                (maintr_rst),
      .UG_maintr_awvalid         (UG_maintr_awvalid),
      .LR_maintr_awready         (LR_maintr_awready),
      .UG_maintr_awaddr          (UG_maintr_awaddr),
      .UG_maintr_wvalid          (UG_maintr_wvalid),
      .LR_maintr_wready          (LR_maintr_wready),
      .UG_maintr_wdata           (UG_maintr_wdata),
      .LR_maintr_bvalid          (LR_maintr_bvalid),
      .UG_maintr_bready          (UG_maintr_bready),
      .LR_maintr_bresp           (LR_maintr_bresp),
      .UG_maintr_arvalid         (UG_maintr_arvalid),
      .LR_maintr_arready         (LR_maintr_arready),
      .UG_maintr_araddr          (UG_maintr_araddr),
      .LR_maintr_rvalid          (LR_maintr_rvalid),
      .UG_maintr_rready          (UG_maintr_rready),
      .LR_maintr_rdata           (LR_maintr_rdata),
      .LR_maintr_rresp           (LR_maintr_rresp),
      .LR_cfgr_awvalid           (LR_cfgr_awvalid),
      .CF_cfgr_awready           (CF_cfgr_awready),
      .LR_cfgr_awaddr            (LR_cfgr_awaddr),
      .LR_cfgr_awprot            (LR_cfgr_awprot),
      .LR_cfgr_wvalid            (LR_cfgr_wvalid),
      .CF_cfgr_wready            (CF_cfgr_wready),
      .LR_cfgr_wdata             (LR_cfgr_wdata),
      .LR_cfgr_wstrb             (LR_cfgr_wstrb),
      .CF_cfgr_bvalid            (CF_cfgr_bvalid),
      .LR_cfgr_bready            (LR_cfgr_bready),
      .CF_cfgr_bresp             (CF_cfgr_bresp),
      .LR_cfgr_arvalid           (LR_cfgr_arvalid),
      .CF_cfgr_arready           (CF_cfgr_arready),
      .LR_cfgr_araddr            (LR_cfgr_araddr),
      .LR_cfgr_arprot            (LR_cfgr_arprot),
      .CF_cfgr_rvalid            (CF_cfgr_rvalid),
      .LR_cfgr_rready            (LR_cfgr_rready),
      .CF_cfgr_rdata             (CF_cfgr_rdata),
      .CF_cfgr_rresp             (CF_cfgr_rresp),
      .LR_lrtx_req_tvalid        (LR_lrtx_req_tvalid),
      .LA_lrtx_req_tready        (LA_lrtx_req_tready),
      .LR_lrtx_req_tdata         (LR_lrtx_req_tdata),
      .LR_lrtx_req_tkeep         (LR_lrtx_req_tkeep),
      .LR_lrtx_req_tlast         (LR_lrtx_req_tlast),
      .LR_lrtx_req_tuser         (LR_lrtx_req_tuser),
      .LR_lrtx_resp_tvalid       (LR_lrtx_resp_tvalid),
      .LA_lrtx_resp_tready       (LA_lrtx_resp_tready),
      .LR_lrtx_resp_tdata        (LR_lrtx_resp_tdata),
      .LR_lrtx_resp_tkeep        (LR_lrtx_resp_tkeep),
      .LR_lrtx_resp_tlast        (LR_lrtx_resp_tlast),
      .LR_lrtx_resp_tuser        (LR_lrtx_resp_tuser),
      .LA_lrrx_tvalid            (LA_lrrx_tvalid),
      .LR_lrrx_tready            (LR_lrrx_tready),
      .LA_lrrx_tdata             (LA_lrrx_tdata),
      .LA_lrrx_tkeep             (LA_lrrx_tkeep),
      .LA_lrrx_tlast             (LA_lrrx_tlast),
      .LA_lrrx_tuser             (LA_lrrx_tuser),
      .LC_deviceid               (LC_deviceid)
     );
   // }}} end log_maint_top instantiation

  // Connect Arbiter ports to log maint ports when maint is enabled
  // TX Request Interface
  //----------------------------------------
  assign UG_tx_portg_tvalid_int  = LR_lrtx_req_tvalid;
  assign LA_lrtx_req_tready      = LA_tx_portg_tready_int;
  assign UG_tx_portg_tdata_int   = LR_lrtx_req_tdata;
  assign UG_tx_portg_tkeep_int   = LR_lrtx_req_tkeep;
  assign UG_tx_portg_tlast_int   = LR_lrtx_req_tlast;
  assign UG_tx_portg_tuser_int   = LR_lrtx_req_tuser;

  // TX Response Interface
  //----------------------------------------
  assign UG_tx_porth_tvalid_int  = LR_lrtx_resp_tvalid;
  assign LA_lrtx_resp_tready     = LA_tx_porth_tready_int;
  assign UG_tx_porth_tdata_int   = LR_lrtx_resp_tdata;
  assign UG_tx_porth_tkeep_int   = LR_lrtx_resp_tkeep;
  assign UG_tx_porth_tlast_int   = LR_lrtx_resp_tlast;
  assign UG_tx_porth_tuser_int   = LR_lrtx_resp_tuser;

  // RX Interface
  //----------------------------------------
  assign LA_lrrx_tvalid          = LA_rx_porth_tvalid_int;
  assign UG_rx_porth_tready_int  = LR_lrrx_tready;
  assign LA_lrrx_tdata           = LA_rx_porth_tdata_int;
  assign LA_lrrx_tkeep           = LA_rx_porth_tkeep_int;
  assign LA_lrrx_tlast           = LA_rx_porth_tlast_int;
  assign LA_lrrx_tuser           = LA_rx_porth_tuser_int;

  // Tie core outputs to 0 when maint is present
  // TX Request Interface
  //----------------------------------------
  assign LA_tx_portg_tready      = 0;

  // TX Response Interface
  //----------------------------------------
  assign LA_tx_porth_tready      = 0;

  // RX Interface
  //----------------------------------------
  assign LA_rx_porth_tvalid      = 0;
  assign LA_rx_porth_tdata       = 0;
  assign LA_rx_porth_tkeep       = 0;
  assign LA_rx_porth_tlast       = 0;
  assign LA_rx_porth_tuser       = 0;

end // end if (MAINT_CFG == 1)
// If the maintenance master block is not enabled from the GUI, do not generate it
else begin: maint_block_disabled_gen // if (MAINT_CFG == 0)

  // Tie off outputs if the maint block is not enabled
  assign LR_maintr_awready = 0;       // Write Port Ready
  assign LR_maintr_wready  = 0;       // Write Port Ready
  assign LR_maintr_bvalid  = 0;       // Write Response Valid
  assign LR_maintr_bresp   = 0;       // Write Response
  assign LR_maintr_arready = 0;       // Read Port Ready
  assign LR_maintr_rvalid  = 0;       // Read Response Valid
  assign LR_maintr_rdata   = 0;       // Read Data
  assign LR_maintr_rresp   = 0;       // Read Response
  assign LR_cfgr_awvalid   = 0;       // Write Command Valid
  assign LR_cfgr_awaddr    = 0;       // Write Address
  assign LR_cfgr_wvalid    = 0;       // Write Data Valid
  assign LR_cfgr_wdata     = 0;       // Write Data
  assign LR_cfgr_wstrb     = 0;       // Write Data byte enables
  assign LR_cfgr_awprot    = 0;       // Write Protection (Tied to 0)
  assign LR_cfgr_bready    = 0;       // Write Response Fabric Ready
  assign LR_cfgr_arvalid   = 0;       // Read Command Valid
  assign LR_cfgr_araddr    = 0;       // Read Address
  assign LR_cfgr_arprot    = 0;       // Read Protection (Tied to 0)
  assign LR_cfgr_rready    = 0;       // Read Response Fabric Ready

  // Connect Arbiter ports to core inputs and outputs when maint is not present
  // TX Request Interface
  //----------------------------------------
  assign UG_tx_portg_tvalid_int  = UG_tx_portg_tvalid;
  assign LA_tx_portg_tready      = LA_tx_portg_tready_int;
  assign UG_tx_portg_tdata_int   = UG_tx_portg_tdata;
  assign UG_tx_portg_tkeep_int   = UG_tx_portg_tkeep;
  assign UG_tx_portg_tlast_int   = UG_tx_portg_tlast;
  assign UG_tx_portg_tuser_int   = UG_tx_portg_tuser;

  // TX Response Interface
  //----------------------------------------
  assign UG_tx_porth_tvalid_int  = UG_tx_porth_tvalid;
  assign LA_tx_porth_tready      = LA_tx_porth_tready_int;
  assign UG_tx_porth_tdata_int   = UG_tx_porth_tdata;
  assign UG_tx_porth_tkeep_int   = UG_tx_porth_tkeep;
  assign UG_tx_porth_tlast_int   = UG_tx_porth_tlast;
  assign UG_tx_porth_tuser_int   = UG_tx_porth_tuser;

  // RX Interface
  //----------------------------------------
  assign LA_rx_porth_tvalid      = LA_rx_porth_tvalid_int;
  assign UG_rx_porth_tready_int  = UG_rx_porth_tready;
  assign LA_rx_porth_tdata       = LA_rx_porth_tdata_int;
  assign LA_rx_porth_tkeep       = LA_rx_porth_tkeep_int;
  assign LA_rx_porth_tlast       = LA_rx_porth_tlast_int;
  assign LA_rx_porth_tuser       = LA_rx_porth_tuser_int;

end endgenerate // end if (MAINT_CFG == 0)

    // {{{ Receive Arbiter Instance ---------
srio_gen2_v4_1_16_arb_rx
  #(
    .TCQ                        (TCQ),

    .DEVICEID_WIDTH             (DEVICEID_WIDTH),
    .RX_PORTA_FALL_THROUGH      (RX_PORTA_FALL_THROUGH),

    .RX_PORTA_ENABLE_FTYPE_SORT (RX_PORTA_ENABLE_FTYPE_SORT),
    .RX_PORTA_FTYPE_SORT1       (RX_PORTA_FTYPE_SORT1),
    .RX_PORTA_FTYPE_SORT2       (RX_PORTA_FTYPE_SORT2),
    .RX_PORTA_FTYPE_SORT3       (RX_PORTA_FTYPE_SORT3),
    .RX_PORTA_FTYPE_SORT4       (RX_PORTA_FTYPE_SORT4),
    .RX_PORTA_FTYPE_SORT5       (RX_PORTA_FTYPE_SORT5),
    .RX_PORTA_FTYPE_SORT6       (RX_PORTA_FTYPE_SORT6),
    .RX_PORTA_FTYPE_SORT7       (RX_PORTA_FTYPE_SORT7),
    .RX_PORTA_ENABLE_TTYPE_SORT (RX_PORTA_ENABLE_TTYPE_SORT),
    .RX_PORTA_TTYPE_SORT1       (RX_PORTA_TTYPE_SORT1),
    .RX_PORTA_TTYPE_SORT2       (RX_PORTA_TTYPE_SORT2),
    .RX_PORTA_TTYPE_SORT3       (RX_PORTA_TTYPE_SORT3),
    .RX_PORTA_TTYPE_SORT4       (RX_PORTA_TTYPE_SORT4),
    .RX_PORTA_TTYPE_SORT5       (RX_PORTA_TTYPE_SORT5),
    .RX_PORTA_TTYPE_SORT6       (RX_PORTA_TTYPE_SORT6),
    .RX_PORTA_TTYPE_SORT7       (RX_PORTA_TTYPE_SORT7),
    .RX_PORTA_ENABLE_STAT_SORT  (RX_PORTA_ENABLE_STAT_SORT),
    .RX_PORTA_STAT_SORT1        (RX_PORTA_STAT_SORT1),
    .RX_PORTA_STAT_SORT2        (RX_PORTA_STAT_SORT2),
    .RX_PORTA_LCSBA_SUPPORT     (RX_PORTA_LCSBA_SUPPORT),

    .RX_PORTB_ENABLE_FTYPE_SORT (RX_PORTB_ENABLE_FTYPE_SORT),
    .RX_PORTB_FTYPE_SORT1       (RX_PORTB_FTYPE_SORT1),
    .RX_PORTB_FTYPE_SORT2       (RX_PORTB_FTYPE_SORT2),
    .RX_PORTB_FTYPE_SORT3       (RX_PORTB_FTYPE_SORT3),
    .RX_PORTB_FTYPE_SORT4       (RX_PORTB_FTYPE_SORT4),
    .RX_PORTB_FTYPE_SORT5       (RX_PORTB_FTYPE_SORT5),
    .RX_PORTB_FTYPE_SORT6       (RX_PORTB_FTYPE_SORT6),
    .RX_PORTB_FTYPE_SORT7       (RX_PORTB_FTYPE_SORT7),
    .RX_PORTB_ENABLE_TTYPE_SORT (RX_PORTB_ENABLE_TTYPE_SORT),
    .RX_PORTB_TTYPE_SORT1       (RX_PORTB_TTYPE_SORT1),
    .RX_PORTB_TTYPE_SORT2       (RX_PORTB_TTYPE_SORT2),
    .RX_PORTB_TTYPE_SORT3       (RX_PORTB_TTYPE_SORT3),
    .RX_PORTB_TTYPE_SORT4       (RX_PORTB_TTYPE_SORT4),
    .RX_PORTB_TTYPE_SORT5       (RX_PORTB_TTYPE_SORT5),
    .RX_PORTB_TTYPE_SORT6       (RX_PORTB_TTYPE_SORT6),
    .RX_PORTB_TTYPE_SORT7       (RX_PORTB_TTYPE_SORT7),
    .RX_PORTB_ENABLE_STAT_SORT  (RX_PORTB_ENABLE_STAT_SORT),
    .RX_PORTB_STAT_SORT1        (RX_PORTB_STAT_SORT1),
    .RX_PORTB_STAT_SORT2        (RX_PORTB_STAT_SORT2),
    .RX_PORTB_LCSBA_SUPPORT     (RX_PORTB_LCSBA_SUPPORT),

    .RX_PORTC_ENABLE_FTYPE_SORT (RX_PORTC_ENABLE_FTYPE_SORT),
    .RX_PORTC_FTYPE_SORT1       (RX_PORTC_FTYPE_SORT1),
    .RX_PORTC_FTYPE_SORT2       (RX_PORTC_FTYPE_SORT2),
    .RX_PORTC_FTYPE_SORT3       (RX_PORTC_FTYPE_SORT3),
    .RX_PORTC_FTYPE_SORT4       (RX_PORTC_FTYPE_SORT4),
    .RX_PORTC_FTYPE_SORT5       (RX_PORTC_FTYPE_SORT5),
    .RX_PORTC_FTYPE_SORT6       (RX_PORTC_FTYPE_SORT6),
    .RX_PORTC_FTYPE_SORT7       (RX_PORTC_FTYPE_SORT7),
    .RX_PORTC_ENABLE_TTYPE_SORT (RX_PORTC_ENABLE_TTYPE_SORT),
    .RX_PORTC_TTYPE_SORT1       (RX_PORTC_TTYPE_SORT1),
    .RX_PORTC_TTYPE_SORT2       (RX_PORTC_TTYPE_SORT2),
    .RX_PORTC_TTYPE_SORT3       (RX_PORTC_TTYPE_SORT3),
    .RX_PORTC_TTYPE_SORT4       (RX_PORTC_TTYPE_SORT4),
    .RX_PORTC_TTYPE_SORT5       (RX_PORTC_TTYPE_SORT5),
    .RX_PORTC_TTYPE_SORT6       (RX_PORTC_TTYPE_SORT6),
    .RX_PORTC_TTYPE_SORT7       (RX_PORTC_TTYPE_SORT7),
    .RX_PORTC_ENABLE_STAT_SORT  (RX_PORTC_ENABLE_STAT_SORT),
    .RX_PORTC_STAT_SORT1        (RX_PORTC_STAT_SORT1),
    .RX_PORTC_STAT_SORT2        (RX_PORTC_STAT_SORT2),
    .RX_PORTC_LCSBA_SUPPORT     (RX_PORTC_LCSBA_SUPPORT),

    .RX_PORTD_ENABLE_FTYPE_SORT (RX_PORTD_ENABLE_FTYPE_SORT),
    .RX_PORTD_FTYPE_SORT1       (RX_PORTD_FTYPE_SORT1),
    .RX_PORTD_FTYPE_SORT2       (RX_PORTD_FTYPE_SORT2),
    .RX_PORTD_FTYPE_SORT3       (RX_PORTD_FTYPE_SORT3),
    .RX_PORTD_FTYPE_SORT4       (RX_PORTD_FTYPE_SORT4),
    .RX_PORTD_FTYPE_SORT5       (RX_PORTD_FTYPE_SORT5),
    .RX_PORTD_FTYPE_SORT6       (RX_PORTD_FTYPE_SORT6),
    .RX_PORTD_FTYPE_SORT7       (RX_PORTD_FTYPE_SORT7),
    .RX_PORTD_ENABLE_TTYPE_SORT (RX_PORTD_ENABLE_TTYPE_SORT),
    .RX_PORTD_TTYPE_SORT1       (RX_PORTD_TTYPE_SORT1),
    .RX_PORTD_TTYPE_SORT2       (RX_PORTD_TTYPE_SORT2),
    .RX_PORTD_TTYPE_SORT3       (RX_PORTD_TTYPE_SORT3),
    .RX_PORTD_TTYPE_SORT4       (RX_PORTD_TTYPE_SORT4),
    .RX_PORTD_TTYPE_SORT5       (RX_PORTD_TTYPE_SORT5),
    .RX_PORTD_TTYPE_SORT6       (RX_PORTD_TTYPE_SORT6),
    .RX_PORTD_TTYPE_SORT7       (RX_PORTD_TTYPE_SORT7),
    .RX_PORTD_ENABLE_STAT_SORT  (RX_PORTD_ENABLE_STAT_SORT),
    .RX_PORTD_STAT_SORT1        (RX_PORTD_STAT_SORT1),
    .RX_PORTD_STAT_SORT2        (RX_PORTD_STAT_SORT2),
    .RX_PORTD_LCSBA_SUPPORT     (RX_PORTD_LCSBA_SUPPORT),

    .RX_PORTE_ENABLE_FTYPE_SORT (RX_PORTE_ENABLE_FTYPE_SORT),
    .RX_PORTE_FTYPE_SORT1       (RX_PORTE_FTYPE_SORT1),
    .RX_PORTE_FTYPE_SORT2       (RX_PORTE_FTYPE_SORT2),
    .RX_PORTE_FTYPE_SORT3       (RX_PORTE_FTYPE_SORT3),
    .RX_PORTE_FTYPE_SORT4       (RX_PORTE_FTYPE_SORT4),
    .RX_PORTE_FTYPE_SORT5       (RX_PORTE_FTYPE_SORT5),
    .RX_PORTE_FTYPE_SORT6       (RX_PORTE_FTYPE_SORT6),
    .RX_PORTE_FTYPE_SORT7       (RX_PORTE_FTYPE_SORT7),
    .RX_PORTE_ENABLE_TTYPE_SORT (RX_PORTE_ENABLE_TTYPE_SORT),
    .RX_PORTE_TTYPE_SORT1       (RX_PORTE_TTYPE_SORT1),
    .RX_PORTE_TTYPE_SORT2       (RX_PORTE_TTYPE_SORT2),
    .RX_PORTE_TTYPE_SORT3       (RX_PORTE_TTYPE_SORT3),
    .RX_PORTE_TTYPE_SORT4       (RX_PORTE_TTYPE_SORT4),
    .RX_PORTE_TTYPE_SORT5       (RX_PORTE_TTYPE_SORT5),
    .RX_PORTE_TTYPE_SORT6       (RX_PORTE_TTYPE_SORT6),
    .RX_PORTE_TTYPE_SORT7       (RX_PORTE_TTYPE_SORT7),
    .RX_PORTE_ENABLE_STAT_SORT  (RX_PORTE_ENABLE_STAT_SORT),
    .RX_PORTE_STAT_SORT1        (RX_PORTE_STAT_SORT1),
    .RX_PORTE_STAT_SORT2        (RX_PORTE_STAT_SORT2),
    .RX_PORTE_LCSBA_SUPPORT     (RX_PORTE_LCSBA_SUPPORT),

    .RX_PORTF_ENABLE_FTYPE_SORT (RX_PORTF_ENABLE_FTYPE_SORT),
    .RX_PORTF_FTYPE_SORT1       (RX_PORTF_FTYPE_SORT1),
    .RX_PORTF_FTYPE_SORT2       (RX_PORTF_FTYPE_SORT2),
    .RX_PORTF_FTYPE_SORT3       (RX_PORTF_FTYPE_SORT3),
    .RX_PORTF_FTYPE_SORT4       (RX_PORTF_FTYPE_SORT4),
    .RX_PORTF_FTYPE_SORT5       (RX_PORTF_FTYPE_SORT5),
    .RX_PORTF_FTYPE_SORT6       (RX_PORTF_FTYPE_SORT6),
    .RX_PORTF_FTYPE_SORT7       (RX_PORTF_FTYPE_SORT7),
    .RX_PORTF_ENABLE_TTYPE_SORT (RX_PORTF_ENABLE_TTYPE_SORT),
    .RX_PORTF_TTYPE_SORT1       (RX_PORTF_TTYPE_SORT1),
    .RX_PORTF_TTYPE_SORT2       (RX_PORTF_TTYPE_SORT2),
    .RX_PORTF_TTYPE_SORT3       (RX_PORTF_TTYPE_SORT3),
    .RX_PORTF_TTYPE_SORT4       (RX_PORTF_TTYPE_SORT4),
    .RX_PORTF_TTYPE_SORT5       (RX_PORTF_TTYPE_SORT5),
    .RX_PORTF_TTYPE_SORT6       (RX_PORTF_TTYPE_SORT6),
    .RX_PORTF_TTYPE_SORT7       (RX_PORTF_TTYPE_SORT7),
    .RX_PORTF_ENABLE_STAT_SORT  (RX_PORTF_ENABLE_STAT_SORT),
    .RX_PORTF_STAT_SORT1        (RX_PORTF_STAT_SORT1),
    .RX_PORTF_STAT_SORT2        (RX_PORTF_STAT_SORT2),
    .RX_PORTF_LCSBA_SUPPORT     (RX_PORTF_LCSBA_SUPPORT),

    .RX_PORTG_ENABLE_FTYPE_SORT (RX_PORTG_ENABLE_FTYPE_SORT),
    .RX_PORTG_FTYPE_SORT1       (RX_PORTG_FTYPE_SORT1),
    .RX_PORTG_FTYPE_SORT2       (RX_PORTG_FTYPE_SORT2),
    .RX_PORTG_FTYPE_SORT3       (RX_PORTG_FTYPE_SORT3),
    .RX_PORTG_FTYPE_SORT4       (RX_PORTG_FTYPE_SORT4),
    .RX_PORTG_FTYPE_SORT5       (RX_PORTG_FTYPE_SORT5),
    .RX_PORTG_FTYPE_SORT6       (RX_PORTG_FTYPE_SORT6),
    .RX_PORTG_FTYPE_SORT7       (RX_PORTG_FTYPE_SORT7),
    .RX_PORTG_ENABLE_TTYPE_SORT (RX_PORTG_ENABLE_TTYPE_SORT),
    .RX_PORTG_TTYPE_SORT1       (RX_PORTG_TTYPE_SORT1),
    .RX_PORTG_TTYPE_SORT2       (RX_PORTG_TTYPE_SORT2),
    .RX_PORTG_TTYPE_SORT3       (RX_PORTG_TTYPE_SORT3),
    .RX_PORTG_TTYPE_SORT4       (RX_PORTG_TTYPE_SORT4),
    .RX_PORTG_TTYPE_SORT5       (RX_PORTG_TTYPE_SORT5),
    .RX_PORTG_TTYPE_SORT6       (RX_PORTG_TTYPE_SORT6),
    .RX_PORTG_TTYPE_SORT7       (RX_PORTG_TTYPE_SORT7),
    .RX_PORTG_ENABLE_STAT_SORT  (RX_PORTG_ENABLE_STAT_SORT),
    .RX_PORTG_STAT_SORT1        (RX_PORTG_STAT_SORT1),
    .RX_PORTG_STAT_SORT2        (RX_PORTG_STAT_SORT2),
    .RX_PORTG_LCSBA_SUPPORT     (RX_PORTG_LCSBA_SUPPORT),

    .RX_PORTH_ENABLE_FTYPE_SORT (RX_PORTH_ENABLE_FTYPE_SORT),
    .RX_PORTH_FTYPE_SORT1       (RX_PORTH_FTYPE_SORT1),
    .RX_PORTH_FTYPE_SORT2       (RX_PORTH_FTYPE_SORT2),
    .RX_PORTH_FTYPE_SORT3       (RX_PORTH_FTYPE_SORT3),
    .RX_PORTH_FTYPE_SORT4       (RX_PORTH_FTYPE_SORT4),
    .RX_PORTH_FTYPE_SORT5       (RX_PORTH_FTYPE_SORT5),
    .RX_PORTH_FTYPE_SORT6       (RX_PORTH_FTYPE_SORT6),
    .RX_PORTH_FTYPE_SORT7       (RX_PORTH_FTYPE_SORT7),
    .RX_PORTH_ENABLE_TTYPE_SORT (RX_PORTH_ENABLE_TTYPE_SORT),
    .RX_PORTH_TTYPE_SORT1       (RX_PORTH_TTYPE_SORT1),
    .RX_PORTH_TTYPE_SORT2       (RX_PORTH_TTYPE_SORT2),
    .RX_PORTH_TTYPE_SORT3       (RX_PORTH_TTYPE_SORT3),
    .RX_PORTH_TTYPE_SORT4       (RX_PORTH_TTYPE_SORT4),
    .RX_PORTH_TTYPE_SORT5       (RX_PORTH_TTYPE_SORT5),
    .RX_PORTH_TTYPE_SORT6       (RX_PORTH_TTYPE_SORT6),
    .RX_PORTH_TTYPE_SORT7       (RX_PORTH_TTYPE_SORT7),
    .RX_PORTH_ENABLE_STAT_SORT  (RX_PORTH_ENABLE_STAT_SORT),
    .RX_PORTH_STAT_SORT1        (RX_PORTH_STAT_SORT1),
    .RX_PORTH_STAT_SORT2        (RX_PORTH_STAT_SORT2),
    .RX_PORTH_LCSBA_SUPPORT     (RX_PORTH_LCSBA_SUPPORT))
  arb_rx_inst
   (
    .log_clk                    (log_clk),
    .log_rst                    (log_rst),

    .LA_rx_porta_tvalid         (LA_rx_porta_tvalid),
    .UG_rx_porta_tready         (UG_rx_porta_tready),
    .LA_rx_porta_tdata          (LA_rx_porta_tdata),
    .LA_rx_porta_tkeep          (LA_rx_porta_tkeep),
    .LA_rx_porta_tlast          (LA_rx_porta_tlast),
    .LA_rx_porta_tuser          (LA_rx_porta_tuser),

    .LA_rx_portb_tvalid         (LA_rx_portb_tvalid),
    .UG_rx_portb_tready         (UG_rx_portb_tready),
    .LA_rx_portb_tdata          (LA_rx_portb_tdata),
    .LA_rx_portb_tkeep          (LA_rx_portb_tkeep),
    .LA_rx_portb_tlast          (LA_rx_portb_tlast),
    .LA_rx_portb_tuser          (LA_rx_portb_tuser),

    .LA_rx_portc_tvalid         (LA_rx_portc_tvalid),
    .UG_rx_portc_tready         (UG_rx_portc_tready),
    .LA_rx_portc_tdata          (LA_rx_portc_tdata),
    .LA_rx_portc_tkeep          (LA_rx_portc_tkeep),
    .LA_rx_portc_tlast          (LA_rx_portc_tlast),
    .LA_rx_portc_tuser          (LA_rx_portc_tuser),

    .LA_rx_portd_tvalid         (LA_rx_portd_tvalid),
    .UG_rx_portd_tready         (UG_rx_portd_tready),
    .LA_rx_portd_tdata          (LA_rx_portd_tdata),
    .LA_rx_portd_tkeep          (LA_rx_portd_tkeep),
    .LA_rx_portd_tlast          (LA_rx_portd_tlast),
    .LA_rx_portd_tuser          (LA_rx_portd_tuser),

    .LA_rx_porte_tvalid         (LA_rx_porte_tvalid),
    .UG_rx_porte_tready         (UG_rx_porte_tready),
    .LA_rx_porte_tdata          (LA_rx_porte_tdata),
    .LA_rx_porte_tkeep          (LA_rx_porte_tkeep),
    .LA_rx_porte_tlast          (LA_rx_porte_tlast),
    .LA_rx_porte_tuser          (LA_rx_porte_tuser),

    .LA_rx_portf_tvalid         (LA_rx_portf_tvalid),
    .UG_rx_portf_tready         (UG_rx_portf_tready),
    .LA_rx_portf_tdata          (LA_rx_portf_tdata),
    .LA_rx_portf_tkeep          (LA_rx_portf_tkeep),
    .LA_rx_portf_tlast          (LA_rx_portf_tlast),
    .LA_rx_portf_tuser          (LA_rx_portf_tuser),

    .LA_rx_portg_tvalid         (LA_rx_portg_tvalid),
    .UG_rx_portg_tready         (UG_rx_portg_tready),
    .LA_rx_portg_tdata          (LA_rx_portg_tdata),
    .LA_rx_portg_tkeep          (LA_rx_portg_tkeep),
    .LA_rx_portg_tlast          (LA_rx_portg_tlast),
    .LA_rx_portg_tuser          (LA_rx_portg_tuser),

    .LA_rx_porth_tvalid         (LA_rx_porth_tvalid_int),
    .UG_rx_porth_tready         (UG_rx_porth_tready_int),
    .LA_rx_porth_tdata          (LA_rx_porth_tdata_int),
    .LA_rx_porth_tkeep          (LA_rx_porth_tkeep_int),
    .LA_rx_porth_tlast          (LA_rx_porth_tlast_int),
    .LA_rx_porth_tuser          (LA_rx_porth_tuser_int),

    .LE_lhrx_tvalid             (LE_lhrx_tvalid),
    .LA_lhrx_tready             (LA_lhrx_tready),
    .LE_lhrx_tdata              (LE_lhrx_tdata),
    .LE_lhrx_tkeep              (LE_lhrx_tkeep),
    .LE_lhrx_tlast              (LE_lhrx_tlast),
    .LE_lhrx_tuser              (LE_lhrx_tuser),
    .LE_unsupported_type        (LE_unsupported_type),

    .LA_port_decode_error       (LA_port_decode_error),

    .LC_lcsba                   (LC_lcsba)
   );
   // }}} ----------------------------------



    // {{{ Transmit Arbiter Instance --------
srio_gen2_v4_1_16_arb_tx
  #(
    .TCQ                     (TCQ),
    .EVAL                    (EVAL),

    .TX_ENABLE_FAIRNESS      (TX_ENABLE_FAIRNESS),// CR# 805160, removed commented code
    //.TX_ENABLE_FAIRNESS      (0), // CR# 805160, commented 

    .TX_PORTA_HELLO          (TX_PORTA_HELLO),
    .TX_PORTB_HELLO          (TX_PORTB_HELLO),
    .TX_PORTC_HELLO          (TX_PORTC_HELLO),
    .TX_PORTD_HELLO          (TX_PORTD_HELLO),
    .TX_PORTE_HELLO          (TX_PORTE_HELLO),
    .TX_PORTF_HELLO          (TX_PORTF_HELLO),
    .TX_PORTG_HELLO          (TX_PORTG_HELLO),
    .TX_PORTH_HELLO          (TX_PORTH_HELLO),

    .TX_PORTA_ENABLE         (TX_PORTA_ENABLE),
    .TX_PORTB_ENABLE         (TX_PORTB_ENABLE),
    .TX_PORTC_ENABLE         (TX_PORTC_ENABLE),
    .TX_PORTD_ENABLE         (TX_PORTD_ENABLE),
    .TX_PORTE_ENABLE         (TX_PORTE_ENABLE),
    .TX_PORTF_ENABLE         (TX_PORTF_ENABLE),
    .TX_PORTG_ENABLE         (TX_PORTG_ENABLE),
    .TX_PORTH_ENABLE         (TX_PORTH_ENABLE),

    .TX_PORTA_PRIORITY       (TX_PORTA_PRIORITY),
    .TX_PORTB_PRIORITY       (TX_PORTB_PRIORITY),
    .TX_PORTC_PRIORITY       (TX_PORTC_PRIORITY),
    .TX_PORTD_PRIORITY       (TX_PORTD_PRIORITY),
    .TX_PORTE_PRIORITY       (TX_PORTE_PRIORITY),
    .TX_PORTF_PRIORITY       (TX_PORTF_PRIORITY),
    .TX_PORTG_PRIORITY       (TX_PORTG_PRIORITY),
    .TX_PORTH_PRIORITY       (TX_PORTH_PRIORITY),

    .TX_PORTA_RESP_CLASS     (TX_PORTA_RESP_CLASS),
    .TX_PORTB_RESP_CLASS     (TX_PORTB_RESP_CLASS),
    .TX_PORTC_RESP_CLASS     (TX_PORTC_RESP_CLASS),
    .TX_PORTD_RESP_CLASS     (TX_PORTD_RESP_CLASS),
    .TX_PORTE_RESP_CLASS     (TX_PORTE_RESP_CLASS),
    .TX_PORTF_RESP_CLASS     (TX_PORTF_RESP_CLASS),
    .TX_PORTG_RESP_CLASS     (TX_PORTG_RESP_CLASS),
    .TX_PORTH_RESP_CLASS     (TX_PORTH_RESP_CLASS),
    .CRF_SUPPORT             (CRF_SUPPORT))

  arb_tx_inst
   (
    .log_clk                 (log_clk),
    .log_rst                 (log_rst),

    .UG_tx_porta_tvalid      (UG_tx_porta_tvalid),
    .LA_tx_porta_tready      (LA_tx_porta_tready),
    .UG_tx_porta_tdata       (UG_tx_porta_tdata),
    .UG_tx_porta_tkeep       (UG_tx_porta_tkeep),
    .UG_tx_porta_tlast       (UG_tx_porta_tlast),
    .UG_tx_porta_tuser       (UG_tx_porta_tuser),

    .UG_tx_portb_tvalid      (UG_tx_portb_tvalid),
    .LA_tx_portb_tready      (LA_tx_portb_tready),
    .UG_tx_portb_tdata       (UG_tx_portb_tdata),
    .UG_tx_portb_tkeep       (UG_tx_portb_tkeep),
    .UG_tx_portb_tlast       (UG_tx_portb_tlast),
    .UG_tx_portb_tuser       (UG_tx_portb_tuser),

    .UG_tx_portc_tvalid      (UG_tx_portc_tvalid),
    .LA_tx_portc_tready      (LA_tx_portc_tready),
    .UG_tx_portc_tdata       (UG_tx_portc_tdata),
    .UG_tx_portc_tkeep       (UG_tx_portc_tkeep),
    .UG_tx_portc_tlast       (UG_tx_portc_tlast),
    .UG_tx_portc_tuser       (UG_tx_portc_tuser),

    .UG_tx_portd_tvalid      (UG_tx_portd_tvalid),
    .LA_tx_portd_tready      (LA_tx_portd_tready),
    .UG_tx_portd_tdata       (UG_tx_portd_tdata),
    .UG_tx_portd_tkeep       (UG_tx_portd_tkeep),
    .UG_tx_portd_tlast       (UG_tx_portd_tlast),
    .UG_tx_portd_tuser       (UG_tx_portd_tuser),

    .UG_tx_porte_tvalid      (UG_tx_porte_tvalid),
    .LA_tx_porte_tready      (LA_tx_porte_tready),
    .UG_tx_porte_tdata       (UG_tx_porte_tdata),
    .UG_tx_porte_tkeep       (UG_tx_porte_tkeep),
    .UG_tx_porte_tlast       (UG_tx_porte_tlast),
    .UG_tx_porte_tuser       (UG_tx_porte_tuser),

    .UG_tx_portf_tvalid      (UG_tx_portf_tvalid),
    .LA_tx_portf_tready      (LA_tx_portf_tready),
    .UG_tx_portf_tdata       (UG_tx_portf_tdata),
    .UG_tx_portf_tkeep       (UG_tx_portf_tkeep),
    .UG_tx_portf_tlast       (UG_tx_portf_tlast),
    .UG_tx_portf_tuser       (UG_tx_portf_tuser),

    .UG_tx_portg_tvalid      (UG_tx_portg_tvalid_int),
    .LA_tx_portg_tready      (LA_tx_portg_tready_int),
    .UG_tx_portg_tdata       (UG_tx_portg_tdata_int),
    .UG_tx_portg_tkeep       (UG_tx_portg_tkeep_int),
    .UG_tx_portg_tlast       (UG_tx_portg_tlast_int),
    .UG_tx_portg_tuser       (UG_tx_portg_tuser_int),

    .UG_tx_porth_tvalid      (UG_tx_porth_tvalid_int),
    .LA_tx_porth_tready      (LA_tx_porth_tready_int),
    .UG_tx_porth_tdata       (UG_tx_porth_tdata_int),
    .UG_tx_porth_tkeep       (UG_tx_porth_tkeep_int),
    .UG_tx_porth_tlast       (UG_tx_porth_tlast_int),
    .UG_tx_porth_tuser       (UG_tx_porth_tuser_int),



    .LA_lhtx_tvalid          (LA_lhtx_tvalid),
    .LD_lhtx_tready          (LD_lhtx_tready),
    .LA_lhtx_tdata           (LA_lhtx_tdata),
    .LA_lhtx_tkeep           (LA_lhtx_tkeep),
    .LA_lhtx_tlast           (LA_lhtx_tlast),
    .LA_lhtx_tuser           (LA_lhtx_tuser),

    .BT_response_only        (BT_response_only),

    .PC_maint_only           (PC_maint_only)
   );
   // }}} ----------------------------------

  // {{{ hello_encoder inst
  //--------------------------------------------
  srio_gen2_v4_1_16_hello_encoder
    #(.TCQ                       (TCQ),
      .DEVICEID_WIDTH            (DEVICEID_WIDTH),
      .TARGET_NREAD              (TARGET_NREAD),
      .TARGET_NWRITE             (TARGET_NWRITE),
      .TARGET_NWRITE_R           (TARGET_NWRITE_R),
      .TARGET_SWRITE             (TARGET_SWRITE),
      .TARGET_DB                 (TARGET_DB),
      .TARGET_DS                 (TARGET_DS),
      .TARGET_ATOMIC             (TARGET_ATOMIC),
      .INIT_NREAD                (INIT_NREAD),
      .INIT_NWRITE_R             (INIT_NWRITE_R),
      .INIT_DB                   (INIT_DB),
      .INIT_ATOMIC               (INIT_ATOMIC),
      .MSG_SINK_SINGLE           (MSG_SINK_SINGLE),
      .MSG_SINK_MULTI            (MSG_SINK_MULTI),
      .MSG_INIT_SINGLE           (MSG_INIT_SINGLE),
      .MSG_INIT_MULTI            (MSG_INIT_MULTI),
      .PORT_IO_HELLO             (PORT_IO_HELLO),
      .PORT_MSG_HELLO            (PORT_MSG_HELLO),
      .PORT_MAINT_HELLO          (PORT_MAINT_HELLO))
    hello_encoder_inst
     (.log_clk                   (log_clk),
      .log_rst                   (log_rst),
      .BR_bufr_tvalid            (BR_bufr_tvalid),
      .LE_bufr_tready            (LE_bufr_tready),
      .BR_bufr_tdata             (BR_bufr_tdata),
      .BR_bufr_tkeep             (BR_bufr_tkeep),
      .BR_bufr_tlast             (BR_bufr_tlast),
      .BR_bufr_tuser             (BR_bufr_tuser),
      .LE_lhrx_tvalid            (LE_lhrx_tvalid),
      .LA_lhrx_tready            (LA_lhrx_tready),
      .LE_lhrx_tdata             (LE_lhrx_tdata),
      .LE_lhrx_tkeep             (LE_lhrx_tkeep),
      .LE_lhrx_tlast             (LE_lhrx_tlast),
      .LE_lhrx_tuser             (LE_lhrx_tuser),
      .LE_unsupported_type       (LE_unsupported_type)
     );
   // }}} end hello_encoder inst

  // {{{ hello_decoder inst
  //--------------------------------------------
  srio_gen2_v4_1_16_hello_decoder
    #(.TCQ                       (TCQ),
      .DEVICEID_WIDTH            (DEVICEID_WIDTH),
      .DECODE_FT02               (DECODE_FT02),
      .DECODE_FT05               (DECODE_FT05),
      .DECODE_FT06               (DECODE_FT06),
      .DECODE_FT08               (DECODE_FT08),
      .DECODE_FT09               (DECODE_FT09),
      .DECODE_FT10               (DECODE_FT10),
      .DECODE_FT11               (DECODE_FT11),
      .DECODE_FT13               (DECODE_FT13),
      .CRF_SUPPORT               (CRF_SUPPORT))// CR# 820838, added the CRF support parameter)
    hello_decoder_inst
     (.log_clk                   (log_clk),
      .log_rst                   (log_rst),
      .LD_buft_tvalid            (LD_buft_tvalid),
      .BT_buft_tready            (BT_buft_tready),
      .LD_buft_tdata             (LD_buft_tdata),
      .LD_buft_tkeep             (LD_buft_tkeep),
      .LD_buft_tlast             (LD_buft_tlast),
      .LD_buft_tuser             (LD_buft_tuser),
      .LA_lhtx_tvalid            (LA_lhtx_tvalid),
      .LD_lhtx_tready            (LD_lhtx_tready),
      .LA_lhtx_tdata             (LA_lhtx_tdata),
      .LA_lhtx_tkeep             (LA_lhtx_tkeep),
      .LA_lhtx_tlast             (LA_lhtx_tlast),
      .LA_lhtx_tuser             (LA_lhtx_tuser)
     );
   // }}} end hello_decoder inst


endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
//
// ARB_TX_MUX
// Description:
// This module uses a mux to arbitrate between ports
//
// Hierarchy:
// LOG_TOP
//    |_____ARB_TX
//             |_____ARB_TX_USER_IF
//             |_____ARB_TX_MUX <-- this module
//    |_____ARB_RX
// ---------------------------------------------------------------------

`timescale 1ps/1ps
// ------------------------------------------------
// below attribute is added to supress the synthesis warnings in vivado tool 8:3332
(* DowngradeIPIdentifiedWarnings="yes" *)
// ------------------------------------------------

module srio_gen2_v4_1_16_arb_tx_mux
  #(
    parameter TCQ                     = 100,  // in pS
    parameter TX_ENABLE_FAIRNESS      = 1,    // when set, use tiebreaking technique {0,1}
    parameter NUMBER_OF_PORTS         = 8)    // total number of ports connected to this module
   (
   // {{{ port declarations ----------------
    // clocks and resets and general signals
    input             log_clk,           // PHY interface clock
    input             log_rst_q,         // Reset for PHY clock Domain

    input             advance_condition, // circumstance that causes the pipeline to move

    // first port object
    input             LAM_port1_tvalid,  // Valid Packet Beat
    input             LAM_port1_tlast,   // Last Beat
    input             LAM_port1_tready,  // Packet Beat Accepted
    input      [3:0]  LAM_port1_id,      // Unique Identifier for each Physical Port

    // second port object
    input             LAM_port2_tvalid,  // Valid Packet Beat
    input             LAM_port2_tlast,   // Last Beat
    input             LAM_port2_tready,  // Packet Beat Accepted
    input      [3:0]  LAM_port2_id,      // Unique Identifier for each Physical Port

    // third port object
    input             LAM_port3_tvalid,  // Valid Packet Beat
    input             LAM_port3_tlast,   // Last Beat
    input             LAM_port3_tready,  // Packet Beat Accepted
    input      [3:0]  LAM_port3_id,      // Unique Identifier for each Physical Port

    // fourth port object
    input             LAM_port4_tvalid,  // Valid Packet Beat
    input             LAM_port4_tlast,   // Last Beat
    input             LAM_port4_tready,  // Packet Beat Accepted
    input      [3:0]  LAM_port4_id,      // Unique Identifier for each Physical Port

    // fifth port object
    input             LAM_port5_tvalid,  // Valid Packet Beat
    input             LAM_port5_tlast,   // Last Beat
    input             LAM_port5_tready,  // Packet Beat Accepted
    input      [3:0]  LAM_port5_id,      // Unique Identifier for each Physical Port

    // sixth port object
    input             LAM_port6_tvalid,  // Valid Packet Beat
    input             LAM_port6_tlast,   // Last Beat
    input             LAM_port6_tready,  // Packet Beat Accepted
    input      [3:0]  LAM_port6_id,      // Unique Identifier for each Physical Port

    // seventh port object
    input             LAM_port7_tvalid,  // Valid Packet Beat
    input             LAM_port7_tlast,   // Last Beat 
    input             LAM_port7_tready,  // Packet Beat Accepted
    input      [3:0]  LAM_port7_id,      // Unique Identifier for each Physical Port

    // eighth port object
    input             LAM_port8_tvalid,  // Valid Packet Beat
    input             LAM_port8_tlast,   // Last Beat
    input             LAM_port8_tready,  // Packet Beat Accepted
    input      [3:0]  LAM_port8_id,      // Unique Identifier for each Physical Port

    output reg [3:0]  LAM_port_winner    // Return Value - holds the Physical Port ID

   // }}} ----------------------------------
   );


  // {{{ local parameters -----------------

  // unique port identifier legend
  localparam PORT1 = 4'h7;
  localparam PORT2 = 4'h6;
  localparam PORT3 = 4'h5;
  localparam PORT4 = 4'h4;
  localparam PORT5 = 4'h3;
  localparam PORT6 = 4'h2;
  localparam PORT7 = 4'h1;
  localparam PORT8 = 4'h0;
  localparam NONE  = 4'hF;

  // }}} End local parameters -------------


  // {{{ wire declarations ----------------

  // holds values of pointers to each port, where tiebreaker1 is the first to
  // win in a tie, while the lowest number tiebreak is the least likely to win.
  reg  [3:0] tiebreaker1_loc;
  reg  [3:0] tiebreaker2_loc;
  reg  [3:0] tiebreaker3_loc;
  reg  [3:0] tiebreaker4_loc;
  reg  [3:0] tiebreaker5_loc;
  reg  [3:0] tiebreaker6_loc;
  reg  [3:0] tiebreaker7_loc;
  reg  [3:0] tiebreaker8_loc;

  reg        tb1_we, tb1_we_d;
  reg        tb2_we, tb2_we_d;
  reg        tb3_we, tb3_we_d;
  reg        tb4_we, tb4_we_d;
  reg        tb5_we, tb5_we_d;
  reg        tb6_we, tb6_we_d;
  reg        tb7_we, tb7_we_d;

  // Winning port pointer
  reg  [3:0] winning_port;
  reg  [3:0] winning_port_q;

  // commonly used signals
  reg        search_for_tvalid;           // When asserted, arbitration begins for next port
  reg        search_for_tvalid_q;         // When asserted, arbitration begins for next port - registered
  reg        find_first_beat;             // used in determining if a packet has begun or not
  reg        out_of_packet;               // asserts when the arbiter is not servicing a packet
  reg        out_of_packet_q;             // asserts when the arbiter is not servicing a packet - registered


  // make a bus of the TVALID and TREADY signals
  wire [7:0] tready_list = {LAM_port1_tready, LAM_port2_tready, LAM_port3_tready, LAM_port4_tready,
                            LAM_port5_tready, LAM_port6_tready, LAM_port7_tready, LAM_port8_tready};
  wire [7:0] tvalid_list = {LAM_port1_tvalid, LAM_port2_tvalid, LAM_port3_tvalid, LAM_port4_tvalid,
                            LAM_port5_tvalid, LAM_port6_tvalid, LAM_port7_tvalid, LAM_port8_tvalid};
  wire [7:0] tlast_list  = {LAM_port1_tlast,  LAM_port2_tlast,  LAM_port3_tlast,  LAM_port4_tlast, 
                            LAM_port5_tlast,  LAM_port6_tlast,  LAM_port7_tlast,  LAM_port8_tlast};

  // }}} End wire declarations ------------


  // {{{ Commonly Used Signal Assignments -

  // indicate when out of packet so we can find the first beat
  always @* begin
    out_of_packet = out_of_packet_q;
    if (tready_list[winning_port] && tlast_list[winning_port] && advance_condition) begin
      out_of_packet = 1'b1;
    end else if (|tvalid_list) begin
      out_of_packet = 1'b0;
    end
  end
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      out_of_packet_q     <= #TCQ 1'b1;
      search_for_tvalid_q <= #TCQ 1'b0;
    end else begin
      out_of_packet_q     <= #TCQ out_of_packet;
      search_for_tvalid_q <= #TCQ search_for_tvalid;
    end
  end
 
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      find_first_beat <= #TCQ 1'b1;
    end else if (find_first_beat && |tvalid_list) begin
      find_first_beat <= #TCQ 1'b0;
    end else if (out_of_packet) begin
      find_first_beat <= #TCQ 1'b1;
    end
  end
 
  // set this when it is ok to start arbitrating for a winning port
// FIXME - CFR probably ok to remove search_for_tvalid
  always @* begin
    search_for_tvalid = search_for_tvalid_q;
    if (!find_first_beat) begin
      search_for_tvalid = 1'b0;
    end else if (|tvalid_list) begin
      search_for_tvalid = 1'b1;
    end
  end

  // }}} End Commonly Used Signals --------


  // {{{ Reorder the tiebreaker -----------
  // reorder tiebreaker list whenever a port gets granted access.
  // winner goes to the back of the list. Each value held within
  // tiebreakerx_loc is a pointer to a port. Each port is assigned
  // to an arbitrary tiebreak location upon reset.
  // In all of the following always blocks, at most, only one 'else if'
  // condition will be implemented. The other option will be removed pre-synth
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      tiebreaker1_loc <= #TCQ PORT1;
    end else if (tb1_we && (NUMBER_OF_PORTS > 1) && (TX_ENABLE_FAIRNESS == 1)) begin
      tiebreaker1_loc <= #TCQ tiebreaker2_loc;
    end
  end

  always @(posedge log_clk) begin
    if (log_rst_q) begin
      tiebreaker2_loc <= #TCQ PORT2;
    end else if (tb2_we && (NUMBER_OF_PORTS > 2) && (TX_ENABLE_FAIRNESS == 1)) begin
      tiebreaker2_loc <= #TCQ tiebreaker3_loc;
    // this condition is only created if this is the final port location
    end else if ((NUMBER_OF_PORTS == 2) && (TX_ENABLE_FAIRNESS == 1)) begin
      casex (tb1_we)
        1'b1     : tiebreaker2_loc <= #TCQ tiebreaker1_loc;
        default  : ;
      endcase
    end
  end

  always @(posedge log_clk) begin
    if (log_rst_q) begin
      tiebreaker3_loc <= #TCQ PORT3;
    end else if (tb3_we && (NUMBER_OF_PORTS > 3) && (TX_ENABLE_FAIRNESS == 1)) begin
      tiebreaker3_loc <= #TCQ tiebreaker4_loc;
    // this condition is only created if this is the final port location
    end else if ((NUMBER_OF_PORTS == 3) && (TX_ENABLE_FAIRNESS == 1)) begin
      casex ({tb1_we, tb2_we})
        2'b1x    : tiebreaker3_loc <= #TCQ tiebreaker1_loc;
        2'b01    : tiebreaker3_loc <= #TCQ tiebreaker2_loc;
        default  : ;
      endcase
    end
  end

  always @(posedge log_clk) begin
    if (log_rst_q) begin
      tiebreaker4_loc <= #TCQ PORT4;
    end else if (tb4_we && (NUMBER_OF_PORTS > 4) && (TX_ENABLE_FAIRNESS == 1)) begin
      tiebreaker4_loc <= #TCQ tiebreaker5_loc;
    // this condition is only created if this is the final port location
    end else if ((NUMBER_OF_PORTS == 4) && (TX_ENABLE_FAIRNESS == 1)) begin
      casex ({tb1_we, tb2_we, tb3_we})
        3'b1xx   : tiebreaker4_loc <= #TCQ tiebreaker1_loc;
        3'b01x   : tiebreaker4_loc <= #TCQ tiebreaker2_loc;
        3'b001   : tiebreaker4_loc <= #TCQ tiebreaker3_loc;
        default  : ;
      endcase
    end
  end

  always @(posedge log_clk) begin
    if (log_rst_q) begin
      tiebreaker5_loc <= #TCQ PORT5;
    end else if (tb5_we && (NUMBER_OF_PORTS > 5) && (TX_ENABLE_FAIRNESS == 1)) begin
      tiebreaker5_loc <= #TCQ tiebreaker6_loc;
    // this condition is only created if this is the final port location
    end else if ((NUMBER_OF_PORTS == 5) && (TX_ENABLE_FAIRNESS == 1)) begin
      casex ({tb1_we, tb2_we, tb3_we, tb4_we})
        4'b1xxx  : tiebreaker5_loc <= #TCQ tiebreaker1_loc;
        4'b01xx  : tiebreaker5_loc <= #TCQ tiebreaker2_loc;
        4'b001x  : tiebreaker5_loc <= #TCQ tiebreaker3_loc;
        4'b0001  : tiebreaker5_loc <= #TCQ tiebreaker4_loc;
        default  : ;
      endcase
    end
  end

  always @(posedge log_clk) begin
    if (log_rst_q) begin
      tiebreaker6_loc <= #TCQ PORT6;
    end else if (tb6_we && (NUMBER_OF_PORTS > 6) && (TX_ENABLE_FAIRNESS == 1)) begin
      tiebreaker6_loc <= #TCQ tiebreaker7_loc;
    // this condition is only created if this is the final port location
    end else if ((NUMBER_OF_PORTS == 6) && (TX_ENABLE_FAIRNESS == 1)) begin
      casex ({tb1_we, tb2_we, tb3_we, tb4_we, tb5_we})
        5'b1xxxx : tiebreaker6_loc <= #TCQ tiebreaker1_loc;
        5'b01xxx : tiebreaker6_loc <= #TCQ tiebreaker2_loc;
        5'b001xx : tiebreaker6_loc <= #TCQ tiebreaker3_loc;
        5'b0001x : tiebreaker6_loc <= #TCQ tiebreaker4_loc;
        5'b00001 : tiebreaker6_loc <= #TCQ tiebreaker5_loc;
        default  : ;
      endcase
    end
  end

  always @(posedge log_clk) begin
    if (log_rst_q) begin
      tiebreaker7_loc <= #TCQ PORT7;
    end else if (tb7_we && (NUMBER_OF_PORTS > 7) && (TX_ENABLE_FAIRNESS == 1)) begin
      tiebreaker7_loc <= #TCQ tiebreaker8_loc;
    // this condition is only created if this is the final port location
    end else if ((NUMBER_OF_PORTS == 7) && (TX_ENABLE_FAIRNESS == 1)) begin
      casex ({tb1_we, tb2_we, tb3_we, tb4_we, tb5_we, tb6_we})
        6'b1xxxxx : tiebreaker7_loc <= #TCQ tiebreaker1_loc;
        6'b01xxxx : tiebreaker7_loc <= #TCQ tiebreaker2_loc;
        6'b001xxx : tiebreaker7_loc <= #TCQ tiebreaker3_loc;
        6'b0001xx : tiebreaker7_loc <= #TCQ tiebreaker4_loc;
        6'b00001x : tiebreaker7_loc <= #TCQ tiebreaker5_loc;
        6'b000001 : tiebreaker7_loc <= #TCQ tiebreaker6_loc;
        default   : ;
      endcase
    end
  end

  always @(posedge log_clk) begin
    if (log_rst_q) begin
      tiebreaker8_loc <= #TCQ PORT8;
    // this condition is only created if this is the final port location
    end else if ((NUMBER_OF_PORTS >= 8) && (TX_ENABLE_FAIRNESS == 1)) begin
      casex ({tb1_we, tb2_we, tb3_we, tb4_we, tb5_we, tb6_we, tb7_we})
        7'b1xxxxxx : tiebreaker8_loc <= #TCQ tiebreaker1_loc;
        7'b01xxxxx : tiebreaker8_loc <= #TCQ tiebreaker2_loc;
        7'b001xxxx : tiebreaker8_loc <= #TCQ tiebreaker3_loc;
        7'b0001xxx : tiebreaker8_loc <= #TCQ tiebreaker4_loc;
        7'b00001xx : tiebreaker8_loc <= #TCQ tiebreaker5_loc;
        7'b000001x : tiebreaker8_loc <= #TCQ tiebreaker6_loc;
        7'b0000001 : tiebreaker8_loc <= #TCQ tiebreaker7_loc;
        default    : ;
      endcase
    end
  end
  // }}} End Reorder the Tiebreaker -------


  // {{{ Set winning_port -----------------
  // find the winning port
  // Any time a higher-numbered port wins, all tiebreakers below
  // it get shifted up. So, set the write enable for all lower ports.
  always @* begin
    winning_port  = winning_port_q;
    tb1_we_d      = 1'b0;
    tb2_we_d      = 1'b0;
    tb3_we_d      = 1'b0;
    tb4_we_d      = 1'b0;
    tb5_we_d      = 1'b0;
    tb6_we_d      = 1'b0;
    tb7_we_d      = 1'b0;
    if (find_first_beat) begin
      if (tvalid_list[tiebreaker1_loc]) begin
        winning_port  = tiebreaker1_loc;
        tb1_we_d      = 1'b1;
        tb2_we_d      = 1'b1;
        tb3_we_d      = 1'b1;
        tb4_we_d      = 1'b1;
        tb5_we_d      = 1'b1;
        tb6_we_d      = 1'b1;
        tb7_we_d      = 1'b1;
      end else if (tvalid_list[tiebreaker2_loc]) begin
        winning_port  = tiebreaker2_loc;
        tb2_we_d      = 1'b1;
        tb3_we_d      = 1'b1;
        tb4_we_d      = 1'b1;
        tb5_we_d      = 1'b1;
        tb6_we_d      = 1'b1;
        tb7_we_d      = 1'b1;
      end else if (tvalid_list[tiebreaker3_loc]) begin
        winning_port  = tiebreaker3_loc;
        tb3_we_d      = 1'b1;
        tb4_we_d      = 1'b1;
        tb5_we_d      = 1'b1;
        tb6_we_d      = 1'b1;
        tb7_we_d      = 1'b1;
      end else if (tvalid_list[tiebreaker4_loc]) begin
        winning_port  = tiebreaker4_loc;
        tb4_we_d      = 1'b1;
        tb5_we_d      = 1'b1;
        tb6_we_d      = 1'b1;
        tb7_we_d      = 1'b1;
      end else if (tvalid_list[tiebreaker5_loc]) begin
        winning_port  = tiebreaker5_loc;
        tb5_we_d      = 1'b1;
        tb6_we_d      = 1'b1;
        tb7_we_d      = 1'b1;
      end else if (tvalid_list[tiebreaker6_loc]) begin
        winning_port  = tiebreaker6_loc;
        tb6_we_d      = 1'b1;
        tb7_we_d      = 1'b1;
      end else if (tvalid_list[tiebreaker7_loc]) begin
        winning_port  = tiebreaker7_loc;
        tb7_we_d      = 1'b1;
      end else begin
//      end else if (tvalid_list[tiebreaker8_loc]) begin
        winning_port  = tiebreaker8_loc;
//      end else begin
//        winning_port  = NONE;
      end
    end
  end
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      //winning_port_q  <= #TCQ NONE;
      winning_port_q  <= #TCQ PORT1;
      tb1_we          <= #TCQ 1'b0;
      tb2_we          <= #TCQ 1'b0;
      tb3_we          <= #TCQ 1'b0;
      tb4_we          <= #TCQ 1'b0;
      tb5_we          <= #TCQ 1'b0;
      tb6_we          <= #TCQ 1'b0;
      tb7_we          <= #TCQ 1'b0;
    end else begin
      winning_port_q  <= #TCQ winning_port;
      tb1_we          <= #TCQ tb1_we_d;
      tb2_we          <= #TCQ tb2_we_d;
      tb3_we          <= #TCQ tb3_we_d;
      tb4_we          <= #TCQ tb4_we_d;
      tb5_we          <= #TCQ tb5_we_d;
      tb6_we          <= #TCQ tb6_we_d;
      tb7_we          <= #TCQ tb7_we_d;
    end
  end

  // Set the winners
  reg [3:0]  lam_port_winner_q;
  always @* begin
    LAM_port_winner = lam_port_winner_q;
    case (winning_port)
      PORT1   : LAM_port_winner = LAM_port1_id;
      PORT2   : LAM_port_winner = LAM_port2_id;
      PORT3   : LAM_port_winner = LAM_port3_id;
      PORT4   : LAM_port_winner = LAM_port4_id;
      PORT5   : LAM_port_winner = LAM_port5_id;
      PORT6   : LAM_port_winner = LAM_port6_id;
      PORT7   : LAM_port_winner = LAM_port7_id;
      //PORT8   : LAM_port_winner = LAM_port8_id;
      default : LAM_port_winner = LAM_port8_id;
      //default : LAM_port_winner = NONE;
    endcase
  end
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      //lam_port_winner_q <= #TCQ NONE;
      lam_port_winner_q <= #TCQ PORT1;
    end else begin
      lam_port_winner_q <= #TCQ LAM_port_winner;
    end
  end

  // }}} End Set winning_port -------------


  // {{{ Coverage and Assertions ----------

    // *- COVERAGE (cg_LAT_tvalid_tiebreaker)
    // Cross all active ports with their location in the tiebreaker list

    // *- COVERAGE (cp_LAT_tiebreak_transition)
    // See a transition from every position to last in the tiebreaker list

    // *- COVERAGE (cp_LAT_higher_tiebreak)
    // Observe a higher tiebreak packet arrive when a lower is already selected

  // }}} End Coverage and Assertions -------------


endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
//
// ARB_TX
// Description:
// This module is strictly used to separate the user from the core.
// It may be replaced by any number of register stages for performance improvement.
//
// Hierarchy:
// LOG_TOP
//    |_____ARB_TX
//             |_____ARB_TX_USER_IF <-- this module
//             |_____ARB_TX_MUX
//    |_____ARB_RX
// ---------------------------------------------------------------------

`timescale 1ps/1ps
// ------------------------------------------------
// below attribute is added to supress the synthesis warnings in vivado tool 8:3332
(* DowngradeIPIdentifiedWarnings="yes" *)
// ------------------------------------------------

module srio_gen2_v4_1_16_arb_tx_user_if
  #(
   // {{{ Parameter declarations -----------
    parameter TCQ                     = 100)  // in pS

   // }}} ----------------------------------
   (
   // {{{ port declarations ----------------
    // clocks and resets and general signals
    input             log_clk,                // PHY interface clock
    input             log_rst_q,              // Reset for PHY clock Domain

    // PORT TX Interface
    input             UG_tx_port_tvalid,      // Valid Packet Beat
    output            LA_tx_port_tready,      // Packet Beat Accepted
    input      [63:0] UG_tx_port_tdata,       // Packet Data
    input       [7:0] UG_tx_port_tkeep,       // Valid bytes in this beat, only valid on last
    input             UG_tx_port_tlast,       // Last Beat
    input      [39:0] UG_tx_port_tuser,       // {DEST_ID, SRC_ID, 5'h0, VC, CRF, 1'b0}

    // 
    input             LA_no_advance,          // hello encoder is stalled
    input             LA_port_mask_tvalid,    // When set, enables tvalid to propigate

    // ARBITER interface
    output reg        UG_tx_port_tvalid_q,    // Valid Packet Beat
    output reg        UG_tx_port_tvalid_raw_q,    // Valid Packet Beat
    input             LA_tx_port_tready_d,    // Packet Beat Accepted
    output reg [63:0] UG_tx_port_tdata_q,     // Packet Data
    output reg  [7:0] UG_tx_port_tkeep_q,     // Valid bytes in this beat, only valid on last
    output reg        UG_tx_port_tlast_q,     // Last Beat
    output reg [39:0] UG_tx_port_tuser_q      // {DEST_ID, SRC_ID, 5'h0, VC, CRF, 1'b0}

   // }}} ----------------------------------
   );


  // {{{ local parameters -----------------

  // }}} End local parameters -------------


  // {{{ wire declarations ----------------
  assign LA_tx_port_tready = (!UG_tx_port_tvalid_raw_q || LA_tx_port_tready_d) && !LA_no_advance; // pull condtion
  wire user_advance_condition =  UG_tx_port_tvalid   && LA_tx_port_tready;   // push condtion
  // }}} End wire declarations ------------

  always @(posedge log_clk) begin
    if (log_rst_q) begin
      UG_tx_port_tvalid_raw_q <= #TCQ 1'b0;
    end else if (user_advance_condition) begin
      UG_tx_port_tvalid_raw_q <= #TCQ 1'b1;
    end else if (LA_tx_port_tready) begin
      UG_tx_port_tvalid_raw_q <= #TCQ 1'b0;
    end
  end
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      UG_tx_port_tvalid_q <= #TCQ 1'b0;
    end else if (user_advance_condition) begin
      UG_tx_port_tvalid_q <= #TCQ LA_port_mask_tvalid;
    end else if (LA_tx_port_tready) begin
      UG_tx_port_tvalid_q <= #TCQ 1'b0;
    end else begin
      UG_tx_port_tvalid_q <= #TCQ UG_tx_port_tvalid_raw_q && LA_port_mask_tvalid;
    end
  end

  always @(posedge log_clk) begin
    if (log_rst_q) begin
      UG_tx_port_tdata_q <= #TCQ 0;
      UG_tx_port_tkeep_q <= #TCQ 0;
      UG_tx_port_tlast_q <= #TCQ 0;
      UG_tx_port_tuser_q <= #TCQ 0;
    end else if (user_advance_condition) begin
      UG_tx_port_tdata_q <= #TCQ UG_tx_port_tdata;
      UG_tx_port_tkeep_q <= #TCQ UG_tx_port_tkeep;
      UG_tx_port_tlast_q <= #TCQ UG_tx_port_tlast;
      UG_tx_port_tuser_q <= #TCQ UG_tx_port_tuser;
    end
  end

endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
//
// ARB_RX
// Description:
// This module holds the transmit logic for the Arbiter
//
// Hierarchy:
// LOG_TOP
//    |_____ARB_TX
//             |_____ARB_TX_USER
//             |_____ARB_TX_MUX
//    |_____ARB_RX <-- this module
// ---------------------------------------------------------------------

`timescale 1ps/1ps

module srio_gen2_v4_1_16_arb_rx
  #(
   // {{{ Parameter declarations -----------
    parameter TCQ                        = 100,        // in pS

    parameter DEVICEID_WIDTH             = 8,          // Source/Destination ID width {8,16}
    parameter RX_PORTA_FALL_THROUGH      = 1,          // If set, all remaining packets fall through to Porta {0,1}

    parameter RX_PORTA_ENABLE_FTYPE_SORT = 7'b1111111, // bitwise enables for ftype search patterns
    parameter RX_PORTA_FTYPE_SORT1       = 1,          // FTYPE search pattern
    parameter RX_PORTA_FTYPE_SORT2       = 1,          // FTYPE search pattern
    parameter RX_PORTA_FTYPE_SORT3       = 1,          // FTYPE search pattern
    parameter RX_PORTA_FTYPE_SORT4       = 1,          // FTYPE search pattern
    parameter RX_PORTA_FTYPE_SORT5       = 1,          // FTYPE search pattern
    parameter RX_PORTA_FTYPE_SORT6       = 1,          // FTYPE search pattern
    parameter RX_PORTA_FTYPE_SORT7       = 1,          // FTYPE search pattern
    parameter RX_PORTA_ENABLE_TTYPE_SORT = 7'b1111111, // bitwise enables for ttype search patterns
    parameter RX_PORTA_TTYPE_SORT1       = 1,          // TTYPE search pattern
    parameter RX_PORTA_TTYPE_SORT2       = 1,          // TTYPE search pattern
    parameter RX_PORTA_TTYPE_SORT3       = 1,          // TTYPE search pattern
    parameter RX_PORTA_TTYPE_SORT4       = 1,          // TTYPE search pattern
    parameter RX_PORTA_TTYPE_SORT5       = 1,          // TTYPE search pattern
    parameter RX_PORTA_TTYPE_SORT6       = 1,          // FTYPE search pattern
    parameter RX_PORTA_TTYPE_SORT7       = 1,          // FTYPE search pattern
    parameter RX_PORTA_ENABLE_STAT_SORT  = 2'b11,      // bitwise enables for stat search patterns
    parameter RX_PORTA_STAT_SORT1        = 1,          // STAT search pattern
    parameter RX_PORTA_STAT_SORT2        = 1,          // STAT search pattern
    parameter RX_PORTA_LCSBA_SUPPORT     = 1,          // If set, I/O can be rerouted to the maint port {0,1}

    parameter RX_PORTB_ENABLE_FTYPE_SORT = 7'b1111111, // bitwise enables for ftype search patterns
    parameter RX_PORTB_FTYPE_SORT1       = 1,          // FTYPE search pattern
    parameter RX_PORTB_FTYPE_SORT2       = 1,          // FTYPE search pattern
    parameter RX_PORTB_FTYPE_SORT3       = 1,          // FTYPE search pattern
    parameter RX_PORTB_FTYPE_SORT4       = 1,          // FTYPE search pattern
    parameter RX_PORTB_FTYPE_SORT5       = 1,          // FTYPE search pattern
    parameter RX_PORTB_FTYPE_SORT6       = 1,          // FTYPE search pattern
    parameter RX_PORTB_FTYPE_SORT7       = 1,          // FTYPE search pattern
    parameter RX_PORTB_ENABLE_TTYPE_SORT = 7'b1111111, // bitwise enables for ttype search patterns
    parameter RX_PORTB_TTYPE_SORT1       = 1,          // TTYPE search pattern
    parameter RX_PORTB_TTYPE_SORT2       = 1,          // TTYPE search pattern
    parameter RX_PORTB_TTYPE_SORT3       = 1,          // TTYPE search pattern
    parameter RX_PORTB_TTYPE_SORT4       = 1,          // TTYPE search pattern
    parameter RX_PORTB_TTYPE_SORT5       = 1,          // TTYPE search pattern
    parameter RX_PORTB_TTYPE_SORT6       = 1,          // TTYPE search pattern
    parameter RX_PORTB_TTYPE_SORT7       = 1,          // TTYPE search pattern
    parameter RX_PORTB_ENABLE_STAT_SORT  = 2'b11,      // bitwise enables for stat search patterns
    parameter RX_PORTB_STAT_SORT1        = 1,          // STAT search pattern
    parameter RX_PORTB_STAT_SORT2        = 1,          // STAT search pattern
    parameter RX_PORTB_LCSBA_SUPPORT     = 1,          // If set, I/O can be rerouted to the maint port {0,1}

    parameter RX_PORTC_ENABLE_FTYPE_SORT = 7'b1111111, // bitwise enables for ftype search patterns
    parameter RX_PORTC_FTYPE_SORT1       = 1,          // FTYPE search pattern
    parameter RX_PORTC_FTYPE_SORT2       = 1,          // FTYPE search pattern
    parameter RX_PORTC_FTYPE_SORT3       = 1,          // FTYPE search pattern
    parameter RX_PORTC_FTYPE_SORT4       = 1,          // FTYPE search pattern
    parameter RX_PORTC_FTYPE_SORT5       = 1,          // FTYPE search pattern
    parameter RX_PORTC_FTYPE_SORT6       = 1,          // FTYPE search pattern
    parameter RX_PORTC_FTYPE_SORT7       = 1,          // FTYPE search pattern
    parameter RX_PORTC_ENABLE_TTYPE_SORT = 7'b1111111, // bitwise enables for ttype search patterns
    parameter RX_PORTC_TTYPE_SORT1       = 1,          // TTYPE search pattern
    parameter RX_PORTC_TTYPE_SORT2       = 1,          // TTYPE search pattern
    parameter RX_PORTC_TTYPE_SORT3       = 1,          // TTYPE search pattern
    parameter RX_PORTC_TTYPE_SORT4       = 1,          // TTYPE search pattern
    parameter RX_PORTC_TTYPE_SORT5       = 1,          // TTYPE search pattern
    parameter RX_PORTC_TTYPE_SORT6       = 1,          // TTYPE search pattern
    parameter RX_PORTC_TTYPE_SORT7       = 1,          // TTYPE search pattern
    parameter RX_PORTC_ENABLE_STAT_SORT  = 2'b11,      // bitwise enables for stat search patterns
    parameter RX_PORTC_STAT_SORT1        = 1,          // STAT search pattern
    parameter RX_PORTC_STAT_SORT2        = 1,          // STAT search pattern
    parameter RX_PORTC_LCSBA_SUPPORT     = 1,          // If set, I/O can be rerouted to the maint port {0,1}

    parameter RX_PORTD_ENABLE_FTYPE_SORT = 7'b1111111, // bitwise enables for ftype search patterns
    parameter RX_PORTD_FTYPE_SORT1       = 1,          // FTYPE search pattern
    parameter RX_PORTD_FTYPE_SORT2       = 1,          // FTYPE search pattern
    parameter RX_PORTD_FTYPE_SORT3       = 1,          // FTYPE search pattern
    parameter RX_PORTD_FTYPE_SORT4       = 1,          // FTYPE search pattern
    parameter RX_PORTD_FTYPE_SORT5       = 1,          // FTYPE search pattern
    parameter RX_PORTD_FTYPE_SORT6       = 1,          // FTYPE search pattern
    parameter RX_PORTD_FTYPE_SORT7       = 1,          // FTYPE search pattern
    parameter RX_PORTD_ENABLE_TTYPE_SORT = 7'b1111111, // bitwise enables for ttype search patterns
    parameter RX_PORTD_TTYPE_SORT1       = 1,          // TTYPE search pattern
    parameter RX_PORTD_TTYPE_SORT2       = 1,          // TTYPE search pattern
    parameter RX_PORTD_TTYPE_SORT3       = 1,          // TTYPE search pattern
    parameter RX_PORTD_TTYPE_SORT4       = 1,          // TTYPE search pattern
    parameter RX_PORTD_TTYPE_SORT5       = 1,          // TTYPE search pattern
    parameter RX_PORTD_TTYPE_SORT6       = 1,          // TTYPE search pattern
    parameter RX_PORTD_TTYPE_SORT7       = 1,          // TTYPE search pattern
    parameter RX_PORTD_ENABLE_STAT_SORT  = 2'b11,      // bitwise enables for stat search patterns
    parameter RX_PORTD_STAT_SORT1        = 1,          // STAT search pattern
    parameter RX_PORTD_STAT_SORT2        = 1,          // STAT search pattern
    parameter RX_PORTD_LCSBA_SUPPORT     = 1,          // If set, I/O can be rerouted to the maint port {0,1}

    parameter RX_PORTE_ENABLE_FTYPE_SORT = 7'b1111111, // bitwise enables for ftype search patterns
    parameter RX_PORTE_FTYPE_SORT1       = 1,          // FTYPE search pattern
    parameter RX_PORTE_FTYPE_SORT2       = 1,          // FTYPE search pattern
    parameter RX_PORTE_FTYPE_SORT3       = 1,          // FTYPE search pattern
    parameter RX_PORTE_FTYPE_SORT4       = 1,          // FTYPE search pattern
    parameter RX_PORTE_FTYPE_SORT5       = 1,          // FTYPE search pattern
    parameter RX_PORTE_FTYPE_SORT6       = 1,          // FTYPE search pattern
    parameter RX_PORTE_FTYPE_SORT7       = 1,          // FTYPE search pattern
    parameter RX_PORTE_ENABLE_TTYPE_SORT = 7'b1111111, // bitwise enables for ttype search patterns
    parameter RX_PORTE_TTYPE_SORT1       = 1,          // TTYPE search pattern
    parameter RX_PORTE_TTYPE_SORT2       = 1,          // TTYPE search pattern
    parameter RX_PORTE_TTYPE_SORT3       = 1,          // TTYPE search pattern
    parameter RX_PORTE_TTYPE_SORT4       = 1,          // TTYPE search pattern
    parameter RX_PORTE_TTYPE_SORT5       = 1,          // TTYPE search pattern
    parameter RX_PORTE_TTYPE_SORT6       = 1,          // TTYPE search pattern
    parameter RX_PORTE_TTYPE_SORT7       = 1,          // TTYPE search pattern
    parameter RX_PORTE_ENABLE_STAT_SORT  = 2'b11,      // bitwise enables for stat search patterns
    parameter RX_PORTE_STAT_SORT1        = 1,          // STAT search pattern
    parameter RX_PORTE_STAT_SORT2        = 1,          // STAT search pattern
    parameter RX_PORTE_LCSBA_SUPPORT     = 1,          // If set, I/O can be rerouted to the maint port {0,1}

    parameter RX_PORTF_ENABLE_FTYPE_SORT = 7'b1111111, // bitwise enables for ftype search patterns
    parameter RX_PORTF_FTYPE_SORT1       = 1,          // FTYPE search pattern
    parameter RX_PORTF_FTYPE_SORT2       = 1,          // FTYPE search pattern
    parameter RX_PORTF_FTYPE_SORT3       = 1,          // FTYPE search pattern
    parameter RX_PORTF_FTYPE_SORT4       = 1,          // FTYPE search pattern
    parameter RX_PORTF_FTYPE_SORT5       = 1,          // FTYPE search pattern
    parameter RX_PORTF_FTYPE_SORT6       = 1,          // FTYPE search pattern
    parameter RX_PORTF_FTYPE_SORT7       = 1,          // FTYPE search pattern
    parameter RX_PORTF_ENABLE_TTYPE_SORT = 7'b1111111, // bitwise enables for ttype search patterns
    parameter RX_PORTF_TTYPE_SORT1       = 1,          // TTYPE search pattern
    parameter RX_PORTF_TTYPE_SORT2       = 1,          // TTYPE search pattern
    parameter RX_PORTF_TTYPE_SORT3       = 1,          // TTYPE search pattern
    parameter RX_PORTF_TTYPE_SORT4       = 1,          // TTYPE search pattern
    parameter RX_PORTF_TTYPE_SORT5       = 1,          // TTYPE search pattern
    parameter RX_PORTF_TTYPE_SORT6       = 1,          // TTYPE search pattern
    parameter RX_PORTF_TTYPE_SORT7       = 1,          // TTYPE search pattern
    parameter RX_PORTF_ENABLE_STAT_SORT  = 2'b11,      // bitwise enables for stat search patterns
    parameter RX_PORTF_STAT_SORT1        = 1,          // STAT search pattern
    parameter RX_PORTF_STAT_SORT2        = 1,          // STAT search pattern
    parameter RX_PORTF_LCSBA_SUPPORT     = 1,          // If set, I/O can be rerouted to the maint port {0,1}

    parameter RX_PORTG_ENABLE_FTYPE_SORT = 7'b1111111, // bitwise enables for ftype search patterns
    parameter RX_PORTG_FTYPE_SORT1       = 1,          // FTYPE search pattern
    parameter RX_PORTG_FTYPE_SORT2       = 1,          // FTYPE search pattern
    parameter RX_PORTG_FTYPE_SORT3       = 1,          // FTYPE search pattern
    parameter RX_PORTG_FTYPE_SORT4       = 1,          // FTYPE search pattern
    parameter RX_PORTG_FTYPE_SORT5       = 1,          // FTYPE search pattern
    parameter RX_PORTG_FTYPE_SORT6       = 1,          // FTYPE search pattern
    parameter RX_PORTG_FTYPE_SORT7       = 1,          // FTYPE search pattern
    parameter RX_PORTG_ENABLE_TTYPE_SORT = 7'b1111111, // bitwise enables for ttype search patterns
    parameter RX_PORTG_TTYPE_SORT1       = 1,          // TTYPE search pattern
    parameter RX_PORTG_TTYPE_SORT2       = 1,          // TTYPE search pattern
    parameter RX_PORTG_TTYPE_SORT3       = 1,          // TTYPE search pattern
    parameter RX_PORTG_TTYPE_SORT4       = 1,          // TTYPE search pattern
    parameter RX_PORTG_TTYPE_SORT5       = 1,          // TTYPE search pattern
    parameter RX_PORTG_TTYPE_SORT6       = 1,          // TTYPE search pattern
    parameter RX_PORTG_TTYPE_SORT7       = 1,          // TTYPE search pattern
    parameter RX_PORTG_ENABLE_STAT_SORT  = 2'b11,      // bitwise enables for stat search patterns
    parameter RX_PORTG_STAT_SORT1        = 1,          // STAT search pattern
    parameter RX_PORTG_STAT_SORT2        = 1,          // STAT search pattern
    parameter RX_PORTG_LCSBA_SUPPORT     = 1,          // If set, I/O can be rerouted to the maint port {0,1}

    parameter RX_PORTH_ENABLE_FTYPE_SORT = 7'b1111111, // bitwise enables for ftype search patterns
    parameter RX_PORTH_FTYPE_SORT1       = 1,          // FTYPE search pattern
    parameter RX_PORTH_FTYPE_SORT2       = 1,          // FTYPE search pattern
    parameter RX_PORTH_FTYPE_SORT3       = 1,          // FTYPE search pattern
    parameter RX_PORTH_FTYPE_SORT4       = 1,          // FTYPE search pattern
    parameter RX_PORTH_FTYPE_SORT5       = 1,          // FTYPE search pattern
    parameter RX_PORTH_FTYPE_SORT6       = 1,          // FTYPE search pattern
    parameter RX_PORTH_FTYPE_SORT7       = 1,          // FTYPE search pattern
    parameter RX_PORTH_ENABLE_TTYPE_SORT = 7'b1111111, // bitwise enables for ttype search patterns
    parameter RX_PORTH_TTYPE_SORT1       = 1,          // TTYPE search pattern
    parameter RX_PORTH_TTYPE_SORT2       = 1,          // TTYPE search pattern
    parameter RX_PORTH_TTYPE_SORT3       = 1,          // TTYPE search pattern
    parameter RX_PORTH_TTYPE_SORT4       = 1,          // TTYPE search pattern
    parameter RX_PORTH_TTYPE_SORT5       = 1,          // TTYPE search pattern
    parameter RX_PORTH_TTYPE_SORT6       = 1,          // TTYPE search pattern
    parameter RX_PORTH_TTYPE_SORT7       = 1,          // TTYPE search pattern
    parameter RX_PORTH_ENABLE_STAT_SORT  = 2'b11,      // bitwise enables for stat search patterns
    parameter RX_PORTH_STAT_SORT1        = 1,          // STAT search pattern
    parameter RX_PORTH_STAT_SORT2        = 1,          // STAT search pattern
    parameter RX_PORTH_LCSBA_SUPPORT     = 1)          // If set, I/O can be rerouted to the maint port {0,1}

   // }}} ----------------------------------
   (
   // {{{ port declarations ----------------
    // clocks and resets and general signals
    input             log_clk,                // PHY interface clock
    input             log_rst,                // Reset for PHY clock Domain

    // PORTA RX Interface
    output reg        LA_rx_porta_tvalid,     // Valid Packet Beat
    input             UG_rx_porta_tready,     // Packet Beat Accepted
    output     [63:0] LA_rx_porta_tdata,      // Packet Data
    output      [7:0] LA_rx_porta_tkeep,      // Valid bytes in this beat, only valid on last
    output reg        LA_rx_porta_tlast,      // Last Beat
    output     [39:0] LA_rx_porta_tuser,      // {DEST_ID, SRC_ID, 5'h0, VC, CRF, 1'b0}

    // PORTB RX Interface
    output reg        LA_rx_portb_tvalid,     // Valid Packet Beat
    input             UG_rx_portb_tready,     // Packet Beat Accepted
    output     [63:0] LA_rx_portb_tdata,      // Packet Data
    output      [7:0] LA_rx_portb_tkeep,      // Valid bytes in this beat, only valid on last
    output reg        LA_rx_portb_tlast,      // Last Beat
    output     [39:0] LA_rx_portb_tuser,      // {DEST_ID, SRC_ID, 5'h0, VC, CRF, 1'b0}

    // PORTC RX Interface
    output reg        LA_rx_portc_tvalid,     // Valid Packet Beat
    input             UG_rx_portc_tready,     // Packet Beat Accepted
    output     [63:0] LA_rx_portc_tdata,      // Packet Data
    output      [7:0] LA_rx_portc_tkeep,      // Valid bytes in this beat, only valid on last
    output reg        LA_rx_portc_tlast,      // Last Beat
    output     [39:0] LA_rx_portc_tuser,      // {DEST_ID, SRC_ID, 5'h0, VC, CRF, 1'b0}

    // PORTD RX Interface
    output reg        LA_rx_portd_tvalid,     // Valid Packet Beat
    input             UG_rx_portd_tready,     // Packet Beat Accepted
    output     [63:0] LA_rx_portd_tdata,      // Packet Data
    output      [7:0] LA_rx_portd_tkeep,      // Valid bytes in this beat, only valid on last
    output reg        LA_rx_portd_tlast,      // Last Beat
    output     [39:0] LA_rx_portd_tuser,      // {DEST_ID, SRC_ID, 5'h0, VC, CRF, 1'b0}

    // PORTE RX Interface
    output reg        LA_rx_porte_tvalid,     // Valid Packet Beat
    input             UG_rx_porte_tready,     // Packet Beat Accepted
    output     [63:0] LA_rx_porte_tdata,      // Packet Data
    output      [7:0] LA_rx_porte_tkeep,      // Valid bytes in this beat, only valid on last
    output reg        LA_rx_porte_tlast,      // Last Beat
    output     [39:0] LA_rx_porte_tuser,      // {DEST_ID, SRC_ID, 5'h0, VC, CRF, 1'b0}

    // PORTF RX Interface
    output reg        LA_rx_portf_tvalid,     // Valid Packet Beat
    input             UG_rx_portf_tready,     // Packet Beat Accepted
    output     [63:0] LA_rx_portf_tdata,      // Packet Data
    output      [7:0] LA_rx_portf_tkeep,      // Valid bytes in this beat, only valid on last
    output reg        LA_rx_portf_tlast,      // Last Beat
    output     [39:0] LA_rx_portf_tuser,      // {DEST_ID, SRC_ID, 5'h0, VC, CRF, 1'b0}

    // PORTG RX Interface
    output reg        LA_rx_portg_tvalid,     // Valid Packet Beat
    input             UG_rx_portg_tready,     // Packet Beat Accepted
    output     [63:0] LA_rx_portg_tdata,      // Packet Data
    output      [7:0] LA_rx_portg_tkeep,      // Valid bytes in this beat, only valid on last
    output reg        LA_rx_portg_tlast,      // Last Beat
    output     [39:0] LA_rx_portg_tuser,      // {DEST_ID, SRC_ID, 5'h0, VC, CRF, 1'b0}

    // PORTH RX Interface
    output reg        LA_rx_porth_tvalid,     // Valid Packet Beat
    input             UG_rx_porth_tready,     // Packet Beat Accepted
    output     [63:0] LA_rx_porth_tdata,      // Packet Data
    output      [7:0] LA_rx_porth_tkeep,      // Valid bytes in this beat, only valid on last
    output reg        LA_rx_porth_tlast,      // Last Beat
    output     [39:0] LA_rx_porth_tuser,      // {DEST_ID, SRC_ID, 5'h0, VC, CRF, 1'b0}


    // Header Encoder RX Interface
    input             LE_lhrx_tvalid,         // Valid Packet Beat
    output            LA_lhrx_tready,         // Packet Beat Accepted
    input      [63:0] LE_lhrx_tdata,          // Packet Data
    input       [7:0] LE_lhrx_tkeep,          // Valid bytes in this beat, only valid on last
    input             LE_lhrx_tlast,          // Last Beat
    input      [39:0] LE_lhrx_tuser,          // {DEST_ID, SRC_ID, 2'h0, HELLO_FMT, 2'h0, VC, CRF, 1'b0}
    input             LE_unsupported_type,    // The packet has been decoded as an unsupported type

    // Error signal
    output reg        LA_port_decode_error,   // No port satisfied the criteria for decode

    input       [9:0] LC_lcsba                // Local Configuration Base Address register mask value

   // }}} ----------------------------------
   );


  // {{{ local parameters -----------------


  // move all of the parameters into an array, to be managed by a generate-for loop
  // parameters can't be two-dimensional. make it flat and bit-select later

  localparam [55:0] RX_PORT_ENABLE_FTYPE_SORT = {RX_PORTH_ENABLE_FTYPE_SORT[6:0], RX_PORTG_ENABLE_FTYPE_SORT[6:0],
                                                 RX_PORTF_ENABLE_FTYPE_SORT[6:0], RX_PORTE_ENABLE_FTYPE_SORT[6:0],
                                                 RX_PORTD_ENABLE_FTYPE_SORT[6:0], RX_PORTC_ENABLE_FTYPE_SORT[6:0],
                                                 RX_PORTB_ENABLE_FTYPE_SORT[6:0], RX_PORTA_ENABLE_FTYPE_SORT[6:0]};

  localparam [31:0] RX_PORT_FTYPE_SORT1 = {RX_PORTH_FTYPE_SORT1[3:0], RX_PORTG_FTYPE_SORT1[3:0],
                                           RX_PORTF_FTYPE_SORT1[3:0], RX_PORTE_FTYPE_SORT1[3:0],
                                           RX_PORTD_FTYPE_SORT1[3:0], RX_PORTC_FTYPE_SORT1[3:0],
                                           RX_PORTB_FTYPE_SORT1[3:0], RX_PORTA_FTYPE_SORT1[3:0]};
  localparam [31:0] RX_PORT_FTYPE_SORT2 = {RX_PORTH_FTYPE_SORT2[3:0], RX_PORTG_FTYPE_SORT2[3:0],
                                           RX_PORTF_FTYPE_SORT2[3:0], RX_PORTE_FTYPE_SORT2[3:0],
                                           RX_PORTD_FTYPE_SORT2[3:0], RX_PORTC_FTYPE_SORT2[3:0],
                                           RX_PORTB_FTYPE_SORT2[3:0], RX_PORTA_FTYPE_SORT2[3:0]};
  localparam [31:0] RX_PORT_FTYPE_SORT3 = {RX_PORTH_FTYPE_SORT3[3:0], RX_PORTG_FTYPE_SORT3[3:0],
                                           RX_PORTF_FTYPE_SORT3[3:0], RX_PORTE_FTYPE_SORT3[3:0],
                                           RX_PORTD_FTYPE_SORT3[3:0], RX_PORTC_FTYPE_SORT3[3:0],
                                           RX_PORTB_FTYPE_SORT3[3:0], RX_PORTA_FTYPE_SORT3[3:0]};
  localparam [31:0] RX_PORT_FTYPE_SORT4 = {RX_PORTH_FTYPE_SORT4[3:0], RX_PORTG_FTYPE_SORT4[3:0],
                                           RX_PORTF_FTYPE_SORT4[3:0], RX_PORTE_FTYPE_SORT4[3:0],
                                           RX_PORTD_FTYPE_SORT4[3:0], RX_PORTC_FTYPE_SORT4[3:0],
                                           RX_PORTB_FTYPE_SORT4[3:0], RX_PORTA_FTYPE_SORT4[3:0]};
  localparam [31:0] RX_PORT_FTYPE_SORT5 = {RX_PORTH_FTYPE_SORT5[3:0], RX_PORTG_FTYPE_SORT5[3:0],
                                           RX_PORTF_FTYPE_SORT5[3:0], RX_PORTE_FTYPE_SORT5[3:0],
                                           RX_PORTD_FTYPE_SORT5[3:0], RX_PORTC_FTYPE_SORT5[3:0],
                                           RX_PORTB_FTYPE_SORT5[3:0], RX_PORTA_FTYPE_SORT5[3:0]};
  localparam [31:0] RX_PORT_FTYPE_SORT6 = {RX_PORTH_FTYPE_SORT6[3:0], RX_PORTG_FTYPE_SORT6[3:0],
                                           RX_PORTF_FTYPE_SORT6[3:0], RX_PORTE_FTYPE_SORT6[3:0],
                                           RX_PORTD_FTYPE_SORT6[3:0], RX_PORTC_FTYPE_SORT6[3:0],
                                           RX_PORTB_FTYPE_SORT6[3:0], RX_PORTA_FTYPE_SORT6[3:0]};
  localparam [31:0] RX_PORT_FTYPE_SORT7 = {RX_PORTH_FTYPE_SORT7[3:0], RX_PORTG_FTYPE_SORT7[3:0],
                                           RX_PORTF_FTYPE_SORT7[3:0], RX_PORTE_FTYPE_SORT7[3:0],
                                           RX_PORTD_FTYPE_SORT7[3:0], RX_PORTC_FTYPE_SORT7[3:0],
                                           RX_PORTB_FTYPE_SORT7[3:0], RX_PORTA_FTYPE_SORT7[3:0]};

  localparam [55:0] RX_PORT_ENABLE_TTYPE_SORT = {RX_PORTH_ENABLE_TTYPE_SORT[6:0], RX_PORTG_ENABLE_TTYPE_SORT[6:0],
                                                 RX_PORTF_ENABLE_TTYPE_SORT[6:0], RX_PORTE_ENABLE_TTYPE_SORT[6:0],
                                                 RX_PORTD_ENABLE_TTYPE_SORT[6:0], RX_PORTC_ENABLE_TTYPE_SORT[6:0],
                                                 RX_PORTB_ENABLE_TTYPE_SORT[6:0], RX_PORTA_ENABLE_TTYPE_SORT[6:0]};

  localparam [31:0] RX_PORT_TTYPE_SORT1 = {RX_PORTH_TTYPE_SORT1[3:0], RX_PORTG_TTYPE_SORT1[3:0],
                                           RX_PORTF_TTYPE_SORT1[3:0], RX_PORTE_TTYPE_SORT1[3:0],
                                           RX_PORTD_TTYPE_SORT1[3:0], RX_PORTC_TTYPE_SORT1[3:0],
                                           RX_PORTB_TTYPE_SORT1[3:0], RX_PORTA_TTYPE_SORT1[3:0]};
  localparam [31:0] RX_PORT_TTYPE_SORT2 = {RX_PORTH_TTYPE_SORT2[3:0], RX_PORTG_TTYPE_SORT2[3:0],
                                           RX_PORTF_TTYPE_SORT2[3:0], RX_PORTE_TTYPE_SORT2[3:0],
                                           RX_PORTD_TTYPE_SORT2[3:0], RX_PORTC_TTYPE_SORT2[3:0],
                                           RX_PORTB_TTYPE_SORT2[3:0], RX_PORTA_TTYPE_SORT2[3:0]};
  localparam [31:0] RX_PORT_TTYPE_SORT3 = {RX_PORTH_TTYPE_SORT3[3:0], RX_PORTG_TTYPE_SORT3[3:0],
                                           RX_PORTF_TTYPE_SORT3[3:0], RX_PORTE_TTYPE_SORT3[3:0],
                                           RX_PORTD_TTYPE_SORT3[3:0], RX_PORTC_TTYPE_SORT3[3:0],
                                           RX_PORTB_TTYPE_SORT3[3:0], RX_PORTA_TTYPE_SORT3[3:0]};
  localparam [31:0] RX_PORT_TTYPE_SORT4 = {RX_PORTH_TTYPE_SORT4[3:0], RX_PORTG_TTYPE_SORT4[3:0],
                                           RX_PORTF_TTYPE_SORT4[3:0], RX_PORTE_TTYPE_SORT4[3:0],
                                           RX_PORTD_TTYPE_SORT4[3:0], RX_PORTC_TTYPE_SORT4[3:0],
                                           RX_PORTB_TTYPE_SORT4[3:0], RX_PORTA_TTYPE_SORT4[3:0]};
  localparam [31:0] RX_PORT_TTYPE_SORT5 = {RX_PORTH_TTYPE_SORT5[3:0], RX_PORTG_TTYPE_SORT5[3:0],
                                           RX_PORTF_TTYPE_SORT5[3:0], RX_PORTE_TTYPE_SORT5[3:0],
                                           RX_PORTD_TTYPE_SORT5[3:0], RX_PORTC_TTYPE_SORT5[3:0],
                                           RX_PORTB_TTYPE_SORT5[3:0], RX_PORTA_TTYPE_SORT5[3:0]};
  localparam [31:0] RX_PORT_TTYPE_SORT6 = {RX_PORTH_TTYPE_SORT6[3:0], RX_PORTG_TTYPE_SORT6[3:0],
                                           RX_PORTF_TTYPE_SORT6[3:0], RX_PORTE_TTYPE_SORT6[3:0],
                                           RX_PORTD_TTYPE_SORT6[3:0], RX_PORTC_TTYPE_SORT6[3:0],
                                           RX_PORTB_TTYPE_SORT6[3:0], RX_PORTA_TTYPE_SORT6[3:0]};
  localparam [31:0] RX_PORT_TTYPE_SORT7 = {RX_PORTH_TTYPE_SORT7[3:0], RX_PORTG_TTYPE_SORT7[3:0],
                                           RX_PORTF_TTYPE_SORT7[3:0], RX_PORTE_TTYPE_SORT7[3:0],
                                           RX_PORTD_TTYPE_SORT7[3:0], RX_PORTC_TTYPE_SORT7[3:0],
                                           RX_PORTB_TTYPE_SORT7[3:0], RX_PORTA_TTYPE_SORT7[3:0]};

  localparam [16:0] RX_PORT_ENABLE_STAT_SORT = {RX_PORTH_ENABLE_STAT_SORT[1:0], RX_PORTG_ENABLE_STAT_SORT[1:0],
                                                RX_PORTF_ENABLE_STAT_SORT[1:0], RX_PORTE_ENABLE_STAT_SORT[1:0],
                                                RX_PORTD_ENABLE_STAT_SORT[1:0], RX_PORTC_ENABLE_STAT_SORT[1:0],
                                                RX_PORTB_ENABLE_STAT_SORT[1:0], RX_PORTA_ENABLE_STAT_SORT[1:0]};

  localparam [31:0] RX_PORT_STAT_SORT1 = {RX_PORTH_STAT_SORT1[3:0], RX_PORTG_STAT_SORT1[3:0],
                                          RX_PORTF_STAT_SORT1[3:0], RX_PORTE_STAT_SORT1[3:0],
                                          RX_PORTD_STAT_SORT1[3:0], RX_PORTC_STAT_SORT1[3:0],
                                          RX_PORTB_STAT_SORT1[3:0], RX_PORTA_STAT_SORT1[3:0]};
  localparam [31:0] RX_PORT_STAT_SORT2 = {RX_PORTH_STAT_SORT2[3:0], RX_PORTG_STAT_SORT2[3:0],
                                          RX_PORTF_STAT_SORT2[3:0], RX_PORTE_STAT_SORT2[3:0],
                                          RX_PORTD_STAT_SORT2[3:0], RX_PORTC_STAT_SORT2[3:0],
                                          RX_PORTB_STAT_SORT2[3:0], RX_PORTA_STAT_SORT2[3:0]};

  localparam [7:0] RX_PORT_FALL_THROUGH = {7'h0, RX_PORTA_FALL_THROUGH[0]};

  localparam [7:0] RX_PORT_LCSBA_SUPPORT = {RX_PORTH_LCSBA_SUPPORT[0], RX_PORTG_LCSBA_SUPPORT[0],
                                            RX_PORTF_LCSBA_SUPPORT[0], RX_PORTE_LCSBA_SUPPORT[0],
                                            RX_PORTD_LCSBA_SUPPORT[0], RX_PORTC_LCSBA_SUPPORT[0],
                                            RX_PORTB_LCSBA_SUPPORT[0], RX_PORTA_LCSBA_SUPPORT[0]};

  // FTYPE declarations
  localparam [3:0] FTYPE_NREAD  = 4'h2;
  localparam [3:0] FTYPE_NWRITE = 4'h5;
  localparam [3:0] FTYPE_DS     = 4'h9;

  // }}} End local parameters -------------


  // {{{ wire declarations ----------------

  reg         log_rst_q = 1;                 // Registered reset signal

  reg  [63:0] le_lhrx_tdata_stg1;            // Registered data
  reg  [39:0] le_lhrx_tuser_stg1;            // Registered user field
  reg   [7:0] le_lhrx_tkeep_stg1;            // Registered strobe
  reg         le_lhrx_tlast_stg1;            // Registered tlast

  reg  [63:0] le_lhrx_tdata_stg2;            // Registered data
  reg  [39:0] le_lhrx_tuser_stg2;            // Registered user field
  reg   [7:0] le_lhrx_tkeep_stg2;            // Registered strobe
  reg         le_lhrx_tlast_stg2;            // Registered tlast

  reg  [63:0] la_rx_portx_tdata;             // final data
  reg  [39:0] la_rx_portx_tuser;             // final user field
  reg   [7:0] la_rx_portx_tkeep;             // final strobe

  wire  [1:0] vacancy_cnt;                   // indicates how many pipeline stages are free
  reg   [1:0] vacancy_cnt_q;                 // indicates how many pipeline stages are free - registered

  wire  [3:0] le_packet_ftype_q;             // Incoming Ftype
  wire  [3:0] le_packet_ttype_q;             // Incoming Ttype
  wire  [3:0] le_packet_stat_q;              // Incoming Stat
  wire [15:0] le_packet_ftype_onehot_q;      // one-hot interpretation of ftype
  wire [15:0] le_packet_ttype_onehot_q;      // one-hot interpretation of ttype
  wire [15:0] le_packet_stat_onehot_q;       // one-hot interpretation of stat
  wire  [9:0] le_packet_lcsba_q;             // Incoming LCSBA
  wire        le_packet_lcsba_hit_q;         // Incoming LCSBA hit
  wire        le_out_of_packet_lhrx_q;       // asserts when the demux is not servicing a packet on lhrx side
  wire        le_find_first_beat_q;          // used in determining if a packet has begun or not

  wire  [7:0] la_rx_port_tvalid_logic_gold;  // array of TVALID determination logic
  wire  [7:0] la_rx_port_tvalid_logic;       // array of TVALID determination logic

  reg         la_rx_porta_tvalid_stg2_d;     // Early version of TVALID - combinatorial
  reg         la_rx_portb_tvalid_stg2_d;     // Early version of TVALID - combinatorial
  reg         la_rx_portc_tvalid_stg2_d;     // Early version of TVALID - combinatorial
  reg         la_rx_portd_tvalid_stg2_d;     // Early version of TVALID - combinatorial
  reg         la_rx_porte_tvalid_stg2_d;     // Early version of TVALID - combinatorial
  reg         la_rx_portf_tvalid_stg2_d;     // Early version of TVALID - combinatorial
  reg         la_rx_portg_tvalid_stg2_d;     // Early version of TVALID - combinatorial
  reg         la_rx_porth_tvalid_stg2_d;     // Early version of TVALID - combinatorial

  reg         la_rx_porta_tvalid_stg2;       // Early version of TVALID
  reg         la_rx_portb_tvalid_stg2;       // Early version of TVALID
  reg         la_rx_portc_tvalid_stg2;       // Early version of TVALID
  reg         la_rx_portd_tvalid_stg2;       // Early version of TVALID
  reg         la_rx_porte_tvalid_stg2;       // Early version of TVALID
  reg         la_rx_portf_tvalid_stg2;       // Early version of TVALID
  reg         la_rx_portg_tvalid_stg2;       // Early version of TVALID
  reg         la_rx_porth_tvalid_stg2;       // Early version of TVALID
  reg         la_rx_port_any_tvalid_stg2;    // any stg2 tvalid is asserted
  reg         la_rx_porta_any_tvalid_stg2;   // any stg2 tvalid is asserted - except porta
  reg         la_rx_portb_any_tvalid_stg2;   // any stg2 tvalid is asserted - except portb
  reg         la_rx_portc_any_tvalid_stg2;   // any stg2 tvalid is asserted - except portc
  reg         la_rx_portd_any_tvalid_stg2;   // any stg2 tvalid is asserted - except portd
  reg         la_rx_porte_any_tvalid_stg2;   // any stg2 tvalid is asserted - except porte
  reg         la_rx_portf_any_tvalid_stg2;   // any stg2 tvalid is asserted - except portf
  reg         la_rx_portg_any_tvalid_stg2;   // any stg2 tvalid is asserted - except portg
  reg         la_rx_porth_any_tvalid_stg2;   // any stg2 tvalid is asserted - except porth

  reg         la_rx_porta_tvalid_stg1_d;     // Early version of TVALID - combinatorial
  reg         la_rx_portb_tvalid_stg1_d;     // Early version of TVALID - combinatorial
  reg         la_rx_portc_tvalid_stg1_d;     // Early version of TVALID - combinatorial
  reg         la_rx_portd_tvalid_stg1_d;     // Early version of TVALID - combinatorial
  reg         la_rx_porte_tvalid_stg1_d;     // Early version of TVALID - combinatorial
  reg         la_rx_portf_tvalid_stg1_d;     // Early version of TVALID - combinatorial
  reg         la_rx_portg_tvalid_stg1_d;     // Early version of TVALID - combinatorial
  reg         la_rx_porth_tvalid_stg1_d;     // Early version of TVALID - combinatorial

  reg         la_rx_porta_tvalid_stg1;       // Early version of TVALID
  reg         la_rx_portb_tvalid_stg1;       // Early version of TVALID
  reg         la_rx_portc_tvalid_stg1;       // Early version of TVALID
  reg         la_rx_portd_tvalid_stg1;       // Early version of TVALID
  reg         la_rx_porte_tvalid_stg1;       // Early version of TVALID
  reg         la_rx_portf_tvalid_stg1;       // Early version of TVALID
  reg         la_rx_portg_tvalid_stg1;       // Early version of TVALID
  reg         la_rx_porth_tvalid_stg1;       // Early version of TVALID
  reg         la_rx_port_any_tvalid_stg1;    // any stg1 tvalid is asserted
  reg         la_rx_porta_any_tvalid_stg1;   // any stg1 tvalid is asserted - except porta
  reg         la_rx_portb_any_tvalid_stg1;   // any stg1 tvalid is asserted - except portb
  reg         la_rx_portc_any_tvalid_stg1;   // any stg1 tvalid is asserted - except portc
  reg         la_rx_portd_any_tvalid_stg1;   // any stg1 tvalid is asserted - except portd
  reg         la_rx_porte_any_tvalid_stg1;   // any stg1 tvalid is asserted - except porte
  reg         la_rx_portf_any_tvalid_stg1;   // any stg1 tvalid is asserted - except portf
  reg         la_rx_portg_any_tvalid_stg1;   // any stg1 tvalid is asserted - except portg
  reg         la_rx_porth_any_tvalid_stg1;   // any stg1 tvalid is asserted - except porth

  wire         la_rx_porta_tvalid_stg0;       // Early version of TVALID
  reg         la_rx_portb_tvalid_stg0;       // Early version of TVALID
  reg         la_rx_portc_tvalid_stg0;       // Early version of TVALID
  wire         la_rx_portd_tvalid_stg0;       // Early version of TVALID
  reg         la_rx_porte_tvalid_stg0;       // Early version of TVALID
  reg         la_rx_portf_tvalid_stg0;       // Early version of TVALID
  reg         la_rx_portg_tvalid_stg0;       // Early version of TVALID
  reg         la_rx_porth_tvalid_stg0;       // Early version of TVALID

  wire        la_rx_porta_tvalid_d;          // Valid Packet Beat - combinatorial
  wire        la_rx_portb_tvalid_d;          // Valid Packet Beat - combinatorial
  wire        la_rx_portc_tvalid_d;          // Valid Packet Beat - combinatorial
  wire        la_rx_portd_tvalid_d;          // Valid Packet Beat - combinatorial
  wire        la_rx_porte_tvalid_d;          // Valid Packet Beat - combinatorial
  wire        la_rx_portf_tvalid_d;          // Valid Packet Beat - combinatorial
  wire        la_rx_portg_tvalid_d;          // Valid Packet Beat - combinatorial
  wire        la_rx_porth_tvalid_d;          // Valid Packet Beat - combinatorial

  wire        la_rx_porta_tlast_d;           // Last Beat - combinatorial
  wire        la_rx_portb_tlast_d;           // Last Beat - combinatorial
  wire        la_rx_portc_tlast_d;           // Last Beat - combinatorial
  wire        la_rx_portd_tlast_d;           // Last Beat - combinatorial
  wire        la_rx_porte_tlast_d;           // Last Beat - combinatorial
  wire        la_rx_portf_tlast_d;           // Last Beat - combinatorial
  wire        la_rx_portg_tlast_d;           // Last Beat - combinatorial
  wire        la_rx_porth_tlast_d;           // Last Beat - combinatorial

  reg         port_decode_error_d;           // detected an error condition
  reg         clear_on_error;                // upon detecting an error, summarily accept the rx packet

  wire        le_lhrx_tvalid_q;
  reg         la_lhrx_tready_d;
  wire [63:0] le_lhrx_tdata_q;
  wire  [7:0] le_lhrx_tkeep_q;
  wire        le_lhrx_tlast_q;
  wire [39:0] le_lhrx_tuser_q;
  wire        le_unsupported_type_q;

  wire        lhrx_advance          = la_lhrx_tready_d && le_lhrx_tvalid_q;
  wire        lhrx_advance_unqual   = la_lhrx_tready_d && le_lhrx_tvalid_q && !port_decode_error_d && !clear_on_error;

  wire  [7:0] tvalid_list = {LA_rx_porta_tvalid, LA_rx_portb_tvalid, LA_rx_portc_tvalid, LA_rx_portd_tvalid,
                             LA_rx_porte_tvalid, LA_rx_portf_tvalid, LA_rx_portg_tvalid, LA_rx_porth_tvalid};
  wire  [7:0] tready_list = {UG_rx_porta_tready, UG_rx_portb_tready, UG_rx_portc_tready, UG_rx_portd_tready,
                             UG_rx_porte_tready, UG_rx_portf_tready, UG_rx_portg_tready, UG_rx_porth_tready};
  wire  [7:0] tlast_list  = {LA_rx_porta_tlast, LA_rx_portb_tlast, LA_rx_portc_tlast, LA_rx_portd_tlast,
                             LA_rx_porte_tlast, LA_rx_portf_tlast, LA_rx_portg_tlast, LA_rx_porth_tlast};

  // }}} End wire declarations ------------


  // {{{ Reset Structure ------------------

  // by rule, we must register the resets before we use them. This is not a
  // synchronizing circuit but rather a method to reduce fanout on the resets.
  always @(posedge log_clk or posedge log_rst) begin
    if (log_rst)
      log_rst_q <= #TCQ 1'b1;
    else
      log_rst_q <= #TCQ 1'b0;
  end

  // }}} End of Reset Structure -----------


  // {{{ Pipeline Instantiation -------------------

  srio_gen2_v4_1_16_arb_rx_pipe
    #(.TCQ                     (TCQ),
      .DEVICEID_WIDTH          (DEVICEID_WIDTH))
    arb_rx_pipe_inst
    (.log_clk                  (log_clk),
     .log_rst_q                (log_rst_q),

     .LC_lcsba                 (LC_lcsba),

     .LE_lhrx_tvalid           (LE_lhrx_tvalid),
     .LA_lhrx_tready           (LA_lhrx_tready),
     .LE_lhrx_tdata            (LE_lhrx_tdata),
     .LE_lhrx_tkeep            (LE_lhrx_tkeep),
     .LE_lhrx_tlast            (LE_lhrx_tlast),
     .LE_lhrx_tuser            (LE_lhrx_tuser),
     .LE_unsupported_type      (LE_unsupported_type),

     .LE_lhrx_tvalid_q         (le_lhrx_tvalid_q),
     .LA_lhrx_tready_d         (la_lhrx_tready_d),
     .LE_lhrx_tdata_q          (le_lhrx_tdata_q),
     .LE_lhrx_tkeep_q          (le_lhrx_tkeep_q),
     .LE_lhrx_tlast_q          (le_lhrx_tlast_q),
     .LE_lhrx_tuser_q          (le_lhrx_tuser_q),
     .LE_unsupported_type_q    (le_unsupported_type_q),

     .LE_packet_ftype_q        (le_packet_ftype_q),
     .LE_packet_ttype_q        (le_packet_ttype_q),
     .LE_packet_stat_q         (le_packet_stat_q),
     .LE_packet_ftype_onehot_q (le_packet_ftype_onehot_q),
     .LE_packet_ttype_onehot_q (le_packet_ttype_onehot_q),
     .LE_packet_stat_onehot_q  (le_packet_stat_onehot_q),
     .LE_packet_lcsba_q        (le_packet_lcsba_q),
     .LE_packet_lcsba_hit_q    (le_packet_lcsba_hit_q),
     .LE_out_of_packet_lhrx_q  (le_out_of_packet_lhrx_q),
     .LE_find_first_beat_q     (le_find_first_beat_q)
   );
  // }}} End of Pipeline Instantiation ------------


  // {{{ Datapath -------------------------

  // the arbiter can store up to two extra beats before it must restrict flow.
  // Data is pushed by the tvalid/tready combination at the source
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      le_lhrx_tdata_stg1 <= #TCQ 0;
      le_lhrx_tuser_stg1 <= #TCQ 0;
      le_lhrx_tkeep_stg1 <= #TCQ 0;
      le_lhrx_tlast_stg1 <= #TCQ 0;

      le_lhrx_tdata_stg2 <= #TCQ 0;
      le_lhrx_tuser_stg2 <= #TCQ 0;
      le_lhrx_tkeep_stg2 <= #TCQ 0;
      le_lhrx_tlast_stg2 <= #TCQ 0;
    end else if (lhrx_advance_unqual) begin
      le_lhrx_tdata_stg1 <= #TCQ le_lhrx_tdata_q;
      le_lhrx_tuser_stg1 <= #TCQ le_lhrx_tuser_q;
      le_lhrx_tkeep_stg1 <= #TCQ le_lhrx_tkeep_q;
      le_lhrx_tlast_stg1 <= #TCQ le_lhrx_tlast_q;

      le_lhrx_tdata_stg2 <= #TCQ le_lhrx_tdata_stg1;
      le_lhrx_tuser_stg2 <= #TCQ le_lhrx_tuser_stg1;
      le_lhrx_tkeep_stg2 <= #TCQ le_lhrx_tkeep_stg1;
      le_lhrx_tlast_stg2 <= #TCQ le_lhrx_tlast_stg1;
    end
  end

  // determine what to present on the outgoing bus(es) based on how many beats are stored.
  // If 0, take directly from the input ports (stage0)
  // If 1, take either stage0 or stage1, depending on the previous value of the vacancy count
  // If 2, take either stage1 or stage2, depending on the previous value of the vacancy count
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      la_rx_portx_tdata  <= #TCQ 64'h0;
      la_rx_portx_tuser  <= #TCQ 40'h0;
      la_rx_portx_tkeep  <= #TCQ 8'h0;
    end else begin
      la_rx_portx_tdata <= #TCQ vacancy_cnt   == 2'h0                          ? la_rx_portx_tdata  :
                                vacancy_cnt   == 2'h1 && vacancy_cnt_q == 2'h0 ? le_lhrx_tdata_q    :
                                vacancy_cnt   == 2'h1 && vacancy_cnt_q != 2'h0 &&
                                !lhrx_advance_unqual                           ? le_lhrx_tdata_stg1 :
                                vacancy_cnt   == 2'h1                          ? le_lhrx_tdata_q    :
                                vacancy_cnt_q == 2'h1                          ? le_lhrx_tdata_stg1 :
                                                                                 le_lhrx_tdata_stg2;
      la_rx_portx_tuser <= #TCQ vacancy_cnt   == 2'h0                          ? la_rx_portx_tuser  :
                                vacancy_cnt   == 2'h1 && vacancy_cnt_q == 2'h0 ? le_lhrx_tuser_q    :
                                vacancy_cnt   == 2'h1 && vacancy_cnt_q != 2'h0 &&
                                !lhrx_advance_unqual                           ? le_lhrx_tuser_stg1 :
                                vacancy_cnt   == 2'h1                          ? le_lhrx_tuser_q    :
                                vacancy_cnt_q == 2'h1                          ? le_lhrx_tuser_stg1 :
                                                                                 le_lhrx_tuser_stg2;
      la_rx_portx_tkeep <= #TCQ vacancy_cnt   == 2'h0                          ? la_rx_portx_tkeep  :
                                vacancy_cnt   == 2'h1 && vacancy_cnt_q == 2'h0 ? le_lhrx_tkeep_q    :
                                vacancy_cnt   == 2'h1 && vacancy_cnt_q != 2'h0 &&
                                !lhrx_advance_unqual                           ? le_lhrx_tkeep_stg1 :
                                vacancy_cnt   == 2'h1                          ? le_lhrx_tkeep_q    :
                                vacancy_cnt_q == 2'h1                          ? le_lhrx_tkeep_stg1 :
                                                                                 le_lhrx_tkeep_stg2;
    end
  end

  // NOTE - if there are timing problems, seperate data into distinct registers
  assign LA_rx_porta_tdata = la_rx_portx_tdata;
  assign LA_rx_portb_tdata = la_rx_portx_tdata;
  assign LA_rx_portc_tdata = la_rx_portx_tdata;
  assign LA_rx_portd_tdata = la_rx_portx_tdata;
  assign LA_rx_porte_tdata = la_rx_portx_tdata;
  assign LA_rx_portf_tdata = la_rx_portx_tdata;
  assign LA_rx_portg_tdata = la_rx_portx_tdata;
  assign LA_rx_porth_tdata = la_rx_portx_tdata;

  assign LA_rx_porta_tuser = la_rx_portx_tuser;
  assign LA_rx_portb_tuser = la_rx_portx_tuser;
  assign LA_rx_portc_tuser = la_rx_portx_tuser;
  assign LA_rx_portd_tuser = la_rx_portx_tuser;
  assign LA_rx_porte_tuser = la_rx_portx_tuser;
  assign LA_rx_portf_tuser = la_rx_portx_tuser;
  assign LA_rx_portg_tuser = la_rx_portx_tuser;
  assign LA_rx_porth_tuser = la_rx_portx_tuser;

  assign LA_rx_porta_tkeep = la_rx_portx_tkeep;
  assign LA_rx_portb_tkeep = la_rx_portx_tkeep;
  assign LA_rx_portc_tkeep = la_rx_portx_tkeep;
  assign LA_rx_portd_tkeep = la_rx_portx_tkeep;
  assign LA_rx_porte_tkeep = la_rx_portx_tkeep;
  assign LA_rx_portf_tkeep = la_rx_portx_tkeep;
  assign LA_rx_portg_tkeep = la_rx_portx_tkeep;
  assign LA_rx_porth_tkeep = la_rx_portx_tkeep;
  // }}} End of Datapath ------------------


  // {{{ Demux Logic ----------------------

  // BIG NASTY COMPARE -
  // repeat the following equation for all eight port decodes:
  // FALL_THROUGH || (FTYPE[ii] && TTYPE[ii] && (STAT[1] || STAT[2])) || LSCBA
  genvar ii;
  generate for (ii = 0; ii < 8; ii = ii+1) begin: demux_decode_gen
    integer ftype_sort1 = RX_PORT_FTYPE_SORT1[ii*4+:4];
    integer ftype_sort2 = RX_PORT_FTYPE_SORT2[ii*4+:4];
    integer ftype_sort3 = RX_PORT_FTYPE_SORT3[ii*4+:4];
    integer ftype_sort4 = RX_PORT_FTYPE_SORT4[ii*4+:4];
    integer ftype_sort5 = RX_PORT_FTYPE_SORT5[ii*4+:4];
    integer ftype_sort6 = RX_PORT_FTYPE_SORT6[ii*4+:4];
    integer ftype_sort7 = RX_PORT_FTYPE_SORT7[ii*4+:4];

    integer ttype_sort1 = RX_PORT_TTYPE_SORT1[ii*4+:4];
    integer ttype_sort2 = RX_PORT_TTYPE_SORT2[ii*4+:4];
    integer ttype_sort3 = RX_PORT_TTYPE_SORT3[ii*4+:4];
    integer ttype_sort4 = RX_PORT_TTYPE_SORT4[ii*4+:4];
    integer ttype_sort5 = RX_PORT_TTYPE_SORT5[ii*4+:4];
    integer ttype_sort6 = RX_PORT_TTYPE_SORT6[ii*4+:4];
    integer ttype_sort7 = RX_PORT_TTYPE_SORT7[ii*4+:4];

    integer stat_sort1 = RX_PORT_STAT_SORT1[ii*4+:4];
    integer stat_sort2 = RX_PORT_STAT_SORT2[ii*4+:4];

    assign la_rx_port_tvalid_logic[ii] = 
      RX_PORT_FALL_THROUGH[ii] ||

      // FTYPE, TTYPE and STAT are coupled together. All must match to be considered a hit.
      // If TTYPE is not a consideration, keep the corresponding ENABLE_TTYPE_SORT value at zero
      // If STAT  is not a consideration, keep the corresponding ENABLE_STAT_SORT  value at zero
      (!le_unsupported_type_q &&
      // *** Logical Equivalent of ***
      // FTYPE_SORT1 && TTYPE_SORT1 && (STAT_SORT1 || STAT_SORT2)
      (((RX_PORT_ENABLE_FTYPE_SORT[ii*7+0] == 1 && le_packet_ftype_onehot_q[ftype_sort1]) &&
        (RX_PORT_ENABLE_TTYPE_SORT[ii*7+0] != 1 || le_packet_ttype_onehot_q[ttype_sort1]) &&
        ((RX_PORT_ENABLE_STAT_SORT[ii*2+0] != 1 || le_packet_stat_onehot_q[stat_sort1])  &&
         (RX_PORT_ENABLE_STAT_SORT[ii*2+1] != 1 || le_packet_stat_onehot_q[stat_sort2]))) ||

      // *** Logical Equivalent of ***
      // FTYPE_SORT2 && TTYPE_SORT2 && (STAT_SORT1 || STAT_SORT2)
       ((RX_PORT_ENABLE_FTYPE_SORT[ii*7+1] == 1 && le_packet_ftype_onehot_q[ftype_sort2]) &&
        (RX_PORT_ENABLE_TTYPE_SORT[ii*7+1] != 1 || le_packet_ttype_onehot_q[ttype_sort2]) &&
        ((RX_PORT_ENABLE_STAT_SORT[ii*2+0] != 1 || le_packet_stat_onehot_q[stat_sort1])  &&
         (RX_PORT_ENABLE_STAT_SORT[ii*2+1] != 1 || le_packet_stat_onehot_q[stat_sort2]))) ||

      // *** Logical Equivalent of ***
      // FTYPE_SORT3 && TTYPE_SORT3 && (STAT_SORT1 || STAT_SORT2)
       ((RX_PORT_ENABLE_FTYPE_SORT[ii*7+2] == 1 && le_packet_ftype_onehot_q[ftype_sort3]) &&
        (RX_PORT_ENABLE_TTYPE_SORT[ii*7+2] != 1 || le_packet_ttype_onehot_q[ttype_sort3]) &&
        ((RX_PORT_ENABLE_STAT_SORT[ii*2+0] != 1 || le_packet_stat_onehot_q[stat_sort1])  &&
         (RX_PORT_ENABLE_STAT_SORT[ii*2+1] != 1 || le_packet_stat_onehot_q[stat_sort2]))) ||

      // *** Logical Equivalent of ***
      // FTYPE_SORT4 && TTYPE_SORT4 && (STAT_SORT1 || STAT_SORT2)
       ((RX_PORT_ENABLE_FTYPE_SORT[ii*7+3] == 1 && le_packet_ftype_onehot_q[ftype_sort4]) &&
        (RX_PORT_ENABLE_TTYPE_SORT[ii*7+3] != 1 || le_packet_ttype_onehot_q[ttype_sort4]) &&
        ((RX_PORT_ENABLE_STAT_SORT[ii*2+0] != 1 || le_packet_stat_onehot_q[stat_sort1])  &&
         (RX_PORT_ENABLE_STAT_SORT[ii*2+1] != 1 || le_packet_stat_onehot_q[stat_sort2]))) ||

      // *** Logical Equivalent of ***
      // FTYPE_SORT5 && TTYPE_SORT5 && (STAT_SORT1 || STAT_SORT2)
       ((RX_PORT_ENABLE_FTYPE_SORT[ii*7+4] == 1 && le_packet_ftype_onehot_q[ftype_sort5]) &&
        (RX_PORT_ENABLE_TTYPE_SORT[ii*7+4] != 1 || le_packet_ttype_onehot_q[ttype_sort5]) &&
        ((RX_PORT_ENABLE_STAT_SORT[ii*2+0] != 1 || le_packet_stat_onehot_q[stat_sort1])  &&
         (RX_PORT_ENABLE_STAT_SORT[ii*2+1] != 1 || le_packet_stat_onehot_q[stat_sort2]))) ||

      // *** Logical Equivalent of ***
      // FTYPE_SORT6 && TTYPE_SORT6 && (STAT_SORT1 || STAT_SORT2)
       ((RX_PORT_ENABLE_FTYPE_SORT[ii*7+5] == 1 && le_packet_ftype_onehot_q[ftype_sort6]) &&
        (RX_PORT_ENABLE_TTYPE_SORT[ii*7+5] != 1 || le_packet_ttype_onehot_q[ttype_sort6]) &&
        ((RX_PORT_ENABLE_STAT_SORT[ii*2+0] != 1 || le_packet_stat_onehot_q[stat_sort1])  &&
         (RX_PORT_ENABLE_STAT_SORT[ii*2+1] != 1 || le_packet_stat_onehot_q[stat_sort2]))) ||

      // *** Logical Equivalent of ***
      // FTYPE_SORT7 && TTYPE_SORT7 && (STAT_SORT1 || STAT_SORT2)
       ((RX_PORT_ENABLE_FTYPE_SORT[ii*7+6] == 1 && le_packet_ftype_onehot_q[ftype_sort7]) &&
        (RX_PORT_ENABLE_TTYPE_SORT[ii*7+6] != 1 || le_packet_ttype_onehot_q[ttype_sort7]) &&
        ((RX_PORT_ENABLE_STAT_SORT[ii*2+0] != 1 || le_packet_stat_onehot_q[stat_sort1])  &&
         (RX_PORT_ENABLE_STAT_SORT[ii*2+1] != 1 || le_packet_stat_onehot_q[stat_sort2]))) ||

       // LCSBA decode
// FIXME CFR - delete this when we're happy that the hit correctly replaces the compare
//       (RX_PORT_LCSBA_SUPPORT[ii] && le_lhrx_tuser_q[5] && LC_lcsba == le_packet_lcsba_q &&
       (RX_PORT_LCSBA_SUPPORT[ii] && le_lhrx_tuser_q[5] && le_packet_lcsba_hit_q &&
        ((le_packet_ftype_onehot_q[FTYPE_NREAD]) || (le_packet_ftype_onehot_q[FTYPE_NWRITE])) )));

  end
  endgenerate

  // combinatorial demux. In the case of multiple hits, the higher letter (starting with H) wins
  // If no hits, the result is an error

reg  la_rx_portd_tvalid_stg0_c;
reg  la_rx_porta_tvalid_stg0_c;

  always @* begin
      la_rx_porth_tvalid_stg0 = 1'b0;
      la_rx_portg_tvalid_stg0 = 1'b0;
      la_rx_portf_tvalid_stg0 = 1'b0;
      la_rx_porte_tvalid_stg0 = 1'b0;
      la_rx_portd_tvalid_stg0_c = 1'b0;
      la_rx_portc_tvalid_stg0 = 1'b0;
      la_rx_portb_tvalid_stg0 = 1'b0;
      la_rx_porta_tvalid_stg0_c = 1'b0;
      port_decode_error_d     = 1'b0;
      casex (la_rx_port_tvalid_logic)
      8'b1xxxxxxx : la_rx_porth_tvalid_stg0 = lhrx_advance;
      8'b01xxxxxx : la_rx_portg_tvalid_stg0 = lhrx_advance;
      8'b001xxxxx : la_rx_portf_tvalid_stg0 = lhrx_advance;
      8'b0001xxxx : la_rx_porte_tvalid_stg0 = lhrx_advance;
      8'b00001xxx : la_rx_portd_tvalid_stg0_c = lhrx_advance;
      8'b000001xx : la_rx_portc_tvalid_stg0 = lhrx_advance;
      8'b0000001x : la_rx_portb_tvalid_stg0 = lhrx_advance;
      8'b00000001 : la_rx_porta_tvalid_stg0_c = lhrx_advance;
      default     : port_decode_error_d     = le_find_first_beat_q && lhrx_advance && !(le_packet_ftype_onehot_q[FTYPE_DS] && !le_unsupported_type_q);

    endcase
  end

assign la_rx_portd_tvalid_stg0 = la_rx_portd_tvalid_stg0_c || (le_packet_ftype_onehot_q[FTYPE_DS] && !le_unsupported_type_q) ;

assign la_rx_porta_tvalid_stg0 = la_rx_porta_tvalid_stg0_c && ! la_rx_portd_tvalid_stg0; 


  // valid stages, correspond to the two storage stages for data
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      la_rx_porth_tvalid_stg1     <= #TCQ 1'b0;
      la_rx_portg_tvalid_stg1     <= #TCQ 1'b0;
      la_rx_portf_tvalid_stg1     <= #TCQ 1'b0;
      la_rx_porte_tvalid_stg1     <= #TCQ 1'b0;
      la_rx_portd_tvalid_stg1     <= #TCQ 1'b0;
      la_rx_portc_tvalid_stg1     <= #TCQ 1'b0;
      la_rx_portb_tvalid_stg1     <= #TCQ 1'b0;
      la_rx_porta_tvalid_stg1     <= #TCQ 1'b0;

      la_rx_porth_tvalid_stg2     <= #TCQ 1'b0;
      la_rx_portg_tvalid_stg2     <= #TCQ 1'b0;
      la_rx_portf_tvalid_stg2     <= #TCQ 1'b0;
      la_rx_porte_tvalid_stg2     <= #TCQ 1'b0;
      la_rx_portd_tvalid_stg2     <= #TCQ 1'b0;
      la_rx_portc_tvalid_stg2     <= #TCQ 1'b0;
      la_rx_portb_tvalid_stg2     <= #TCQ 1'b0;
      la_rx_porta_tvalid_stg2     <= #TCQ 1'b0;

      la_rx_port_any_tvalid_stg1  <= #TCQ 1'b0;
      la_rx_porta_any_tvalid_stg1 <= #TCQ 1'b0;
      la_rx_portb_any_tvalid_stg1 <= #TCQ 1'b0;
      la_rx_portc_any_tvalid_stg1 <= #TCQ 1'b0;
      la_rx_portd_any_tvalid_stg1 <= #TCQ 1'b0;
      la_rx_porte_any_tvalid_stg1 <= #TCQ 1'b0;
      la_rx_portf_any_tvalid_stg1 <= #TCQ 1'b0;
      la_rx_portg_any_tvalid_stg1 <= #TCQ 1'b0;
      la_rx_porth_any_tvalid_stg1 <= #TCQ 1'b0;

      la_rx_port_any_tvalid_stg2  <= #TCQ 1'b0;
      la_rx_porta_any_tvalid_stg2 <= #TCQ 1'b0;
      la_rx_portb_any_tvalid_stg2 <= #TCQ 1'b0;
      la_rx_portc_any_tvalid_stg2 <= #TCQ 1'b0;
      la_rx_portd_any_tvalid_stg2 <= #TCQ 1'b0;
      la_rx_porte_any_tvalid_stg2 <= #TCQ 1'b0;
      la_rx_portf_any_tvalid_stg2 <= #TCQ 1'b0;
      la_rx_portg_any_tvalid_stg2 <= #TCQ 1'b0;
      la_rx_porth_any_tvalid_stg2 <= #TCQ 1'b0;
    end else begin
      la_rx_porth_tvalid_stg1     <= #TCQ la_rx_porth_tvalid_stg1_d;
      la_rx_portg_tvalid_stg1     <= #TCQ la_rx_portg_tvalid_stg1_d;
      la_rx_portf_tvalid_stg1     <= #TCQ la_rx_portf_tvalid_stg1_d;
      la_rx_porte_tvalid_stg1     <= #TCQ la_rx_porte_tvalid_stg1_d;
      la_rx_portd_tvalid_stg1     <= #TCQ la_rx_portd_tvalid_stg1_d;
      la_rx_portc_tvalid_stg1     <= #TCQ la_rx_portc_tvalid_stg1_d;
      la_rx_portb_tvalid_stg1     <= #TCQ la_rx_portb_tvalid_stg1_d;
      la_rx_porta_tvalid_stg1     <= #TCQ la_rx_porta_tvalid_stg1_d;

      la_rx_porth_tvalid_stg2     <= #TCQ la_rx_porth_tvalid_stg2_d;
      la_rx_portg_tvalid_stg2     <= #TCQ la_rx_portg_tvalid_stg2_d;
      la_rx_portf_tvalid_stg2     <= #TCQ la_rx_portf_tvalid_stg2_d;
      la_rx_porte_tvalid_stg2     <= #TCQ la_rx_porte_tvalid_stg2_d;
      la_rx_portd_tvalid_stg2     <= #TCQ la_rx_portd_tvalid_stg2_d;
      la_rx_portc_tvalid_stg2     <= #TCQ la_rx_portc_tvalid_stg2_d;
      la_rx_portb_tvalid_stg2     <= #TCQ la_rx_portb_tvalid_stg2_d;
      la_rx_porta_tvalid_stg2     <= #TCQ la_rx_porta_tvalid_stg2_d;

      la_rx_port_any_tvalid_stg1  <= #TCQ (la_rx_porta_tvalid_stg1_d || la_rx_portb_tvalid_stg1_d ||
                                           la_rx_portc_tvalid_stg1_d || la_rx_portd_tvalid_stg1_d ||
                                           la_rx_porte_tvalid_stg1_d || la_rx_portf_tvalid_stg1_d ||
                                           la_rx_portg_tvalid_stg1_d || la_rx_porth_tvalid_stg1_d);
      la_rx_porta_any_tvalid_stg1 <= #TCQ (la_rx_portb_tvalid_stg1_d ||
                                           la_rx_portc_tvalid_stg1_d || la_rx_portd_tvalid_stg1_d ||
                                           la_rx_porte_tvalid_stg1_d || la_rx_portf_tvalid_stg1_d ||
                                           la_rx_portg_tvalid_stg1_d || la_rx_porth_tvalid_stg1_d);
      la_rx_portb_any_tvalid_stg1 <= #TCQ (la_rx_porta_tvalid_stg1_d ||
                                           la_rx_portc_tvalid_stg1_d || la_rx_portd_tvalid_stg1_d ||
                                           la_rx_porte_tvalid_stg1_d || la_rx_portf_tvalid_stg1_d ||
                                           la_rx_portg_tvalid_stg1_d || la_rx_porth_tvalid_stg1_d);
      la_rx_portc_any_tvalid_stg1 <= #TCQ (la_rx_porta_tvalid_stg1_d || la_rx_portb_tvalid_stg1_d ||
                                           la_rx_portd_tvalid_stg1_d ||
                                           la_rx_porte_tvalid_stg1_d || la_rx_portf_tvalid_stg1_d ||
                                           la_rx_portg_tvalid_stg1_d || la_rx_porth_tvalid_stg1_d);
      la_rx_portd_any_tvalid_stg1 <= #TCQ (la_rx_porta_tvalid_stg1_d || la_rx_portb_tvalid_stg1_d ||
                                           la_rx_portc_tvalid_stg1_d ||
                                           la_rx_porte_tvalid_stg1_d || la_rx_portf_tvalid_stg1_d ||
                                           la_rx_portg_tvalid_stg1_d || la_rx_porth_tvalid_stg1_d);
      la_rx_porte_any_tvalid_stg1 <= #TCQ (la_rx_porta_tvalid_stg1_d || la_rx_portb_tvalid_stg1_d ||
                                           la_rx_portc_tvalid_stg1_d || la_rx_portd_tvalid_stg1_d ||
                                           la_rx_portf_tvalid_stg1_d ||
                                           la_rx_portg_tvalid_stg1_d || la_rx_porth_tvalid_stg1_d);
      la_rx_portf_any_tvalid_stg1 <= #TCQ (la_rx_porta_tvalid_stg1_d || la_rx_portb_tvalid_stg1_d ||
                                           la_rx_portc_tvalid_stg1_d || la_rx_portd_tvalid_stg1_d ||
                                           la_rx_porte_tvalid_stg1_d ||
                                           la_rx_portg_tvalid_stg1_d || la_rx_porth_tvalid_stg1_d);
      la_rx_portg_any_tvalid_stg1 <= #TCQ (la_rx_porta_tvalid_stg1_d || la_rx_portb_tvalid_stg1_d ||
                                           la_rx_portc_tvalid_stg1_d || la_rx_portd_tvalid_stg1_d ||
                                           la_rx_porte_tvalid_stg1_d || la_rx_portf_tvalid_stg1_d ||
                                           la_rx_porth_tvalid_stg1_d);
      la_rx_porth_any_tvalid_stg1 <= #TCQ (la_rx_porta_tvalid_stg1_d || la_rx_portb_tvalid_stg1_d ||
                                           la_rx_portc_tvalid_stg1_d || la_rx_portd_tvalid_stg1_d ||
                                           la_rx_porte_tvalid_stg1_d || la_rx_portf_tvalid_stg1_d ||
                                           la_rx_portg_tvalid_stg1_d);

      la_rx_port_any_tvalid_stg2  <= #TCQ (la_rx_porta_tvalid_stg2_d || la_rx_portb_tvalid_stg2_d ||
                                           la_rx_portc_tvalid_stg2_d || la_rx_portd_tvalid_stg2_d ||
                                           la_rx_porte_tvalid_stg2_d || la_rx_portf_tvalid_stg2_d ||
                                           la_rx_portg_tvalid_stg2_d || la_rx_porth_tvalid_stg2_d);
      la_rx_porta_any_tvalid_stg2 <= #TCQ (la_rx_portb_tvalid_stg2_d ||
                                           la_rx_portc_tvalid_stg2_d || la_rx_portd_tvalid_stg2_d ||
                                           la_rx_porte_tvalid_stg2_d || la_rx_portf_tvalid_stg2_d ||
                                           la_rx_portg_tvalid_stg2_d || la_rx_porth_tvalid_stg2_d);
      la_rx_portb_any_tvalid_stg2 <= #TCQ (la_rx_porta_tvalid_stg2_d ||
                                           la_rx_portc_tvalid_stg2_d || la_rx_portd_tvalid_stg2_d ||
                                           la_rx_porte_tvalid_stg2_d || la_rx_portf_tvalid_stg2_d ||
                                           la_rx_portg_tvalid_stg2_d || la_rx_porth_tvalid_stg2_d);
      la_rx_portc_any_tvalid_stg2 <= #TCQ (la_rx_porta_tvalid_stg2_d || la_rx_portb_tvalid_stg2_d ||
                                           la_rx_portd_tvalid_stg2_d ||
                                           la_rx_porte_tvalid_stg2_d || la_rx_portf_tvalid_stg2_d ||
                                           la_rx_portg_tvalid_stg2_d || la_rx_porth_tvalid_stg2_d);
      la_rx_portd_any_tvalid_stg2 <= #TCQ (la_rx_porta_tvalid_stg2_d || la_rx_portb_tvalid_stg2_d ||
                                           la_rx_portc_tvalid_stg2_d ||
                                           la_rx_porte_tvalid_stg2_d || la_rx_portf_tvalid_stg2_d ||
                                           la_rx_portg_tvalid_stg2_d || la_rx_porth_tvalid_stg2_d);
      la_rx_porte_any_tvalid_stg2 <= #TCQ (la_rx_porta_tvalid_stg2_d || la_rx_portb_tvalid_stg2_d ||
                                           la_rx_portc_tvalid_stg2_d || la_rx_portd_tvalid_stg2_d ||
                                           la_rx_portf_tvalid_stg2_d ||
                                           la_rx_portg_tvalid_stg2_d || la_rx_porth_tvalid_stg2_d);
      la_rx_portf_any_tvalid_stg2 <= #TCQ (la_rx_porta_tvalid_stg2_d || la_rx_portb_tvalid_stg2_d ||
                                           la_rx_portc_tvalid_stg2_d || la_rx_portd_tvalid_stg2_d ||
                                           la_rx_porte_tvalid_stg2_d ||
                                           la_rx_portg_tvalid_stg2_d || la_rx_porth_tvalid_stg2_d);
      la_rx_portg_any_tvalid_stg2 <= #TCQ (la_rx_porta_tvalid_stg2_d || la_rx_portb_tvalid_stg2_d ||
                                           la_rx_portc_tvalid_stg2_d || la_rx_portd_tvalid_stg2_d ||
                                           la_rx_porte_tvalid_stg2_d || la_rx_portf_tvalid_stg2_d ||
                                           la_rx_porth_tvalid_stg2_d);
      la_rx_porth_any_tvalid_stg2 <= #TCQ (la_rx_porta_tvalid_stg2_d || la_rx_portb_tvalid_stg2_d ||
                                           la_rx_portc_tvalid_stg2_d || la_rx_portd_tvalid_stg2_d ||
                                           la_rx_porte_tvalid_stg2_d || la_rx_portf_tvalid_stg2_d ||
                                           la_rx_portg_tvalid_stg2_d);
    end
  end

  always @* begin
    if (lhrx_advance_unqual) begin
      // Stage 1
      la_rx_porth_tvalid_stg1_d = la_rx_porth_tvalid_stg0;
      la_rx_portg_tvalid_stg1_d = la_rx_portg_tvalid_stg0;
      la_rx_portf_tvalid_stg1_d = la_rx_portf_tvalid_stg0;
      la_rx_porte_tvalid_stg1_d = la_rx_porte_tvalid_stg0;
      la_rx_portd_tvalid_stg1_d = la_rx_portd_tvalid_stg0;
      la_rx_portc_tvalid_stg1_d = la_rx_portc_tvalid_stg0;
      la_rx_portb_tvalid_stg1_d = la_rx_portb_tvalid_stg0;
      la_rx_porta_tvalid_stg1_d = la_rx_porta_tvalid_stg0;

      // Stage 2 (contains both set and clear logic)
      la_rx_porth_tvalid_stg2_d = la_rx_porth_tvalid_stg1 &&
                                  !(LA_rx_porth_tvalid && UG_rx_porth_tready && vacancy_cnt_q == 2'h1);
      la_rx_portg_tvalid_stg2_d = la_rx_portg_tvalid_stg1 &&
                                  !(LA_rx_portg_tvalid && UG_rx_portg_tready && vacancy_cnt_q == 2'h1);
      la_rx_portf_tvalid_stg2_d = la_rx_portf_tvalid_stg1 &&
                                  !(LA_rx_portf_tvalid && UG_rx_portf_tready && vacancy_cnt_q == 2'h1);
      la_rx_porte_tvalid_stg2_d = la_rx_porte_tvalid_stg1 &&
                                  !(LA_rx_porte_tvalid && UG_rx_porte_tready && vacancy_cnt_q == 2'h1);
      la_rx_portd_tvalid_stg2_d = la_rx_portd_tvalid_stg1 &&
                                  !(LA_rx_portd_tvalid && UG_rx_portd_tready && vacancy_cnt_q == 2'h1);
      la_rx_portc_tvalid_stg2_d = la_rx_portc_tvalid_stg1 &&
                                  !(LA_rx_portc_tvalid && UG_rx_portc_tready && vacancy_cnt_q == 2'h1);
      la_rx_portb_tvalid_stg2_d = la_rx_portb_tvalid_stg1 &&
                                  !(LA_rx_portb_tvalid && UG_rx_portb_tready && vacancy_cnt_q == 2'h1);
      la_rx_porta_tvalid_stg2_d = la_rx_porta_tvalid_stg1 &&
                                  !(LA_rx_porta_tvalid && UG_rx_porta_tready && vacancy_cnt_q == 2'h1);
    // clear the ready if that beat has been successfully sent
    end else begin
      // Stage 1 (contains both set and clear logic)
      la_rx_porth_tvalid_stg1_d = la_rx_porth_tvalid_stg1 &&
                                  !(LA_rx_porth_tvalid && UG_rx_porth_tready && vacancy_cnt_q == 2'h1);
      la_rx_portg_tvalid_stg1_d = la_rx_portg_tvalid_stg1 &&
                                  !(LA_rx_portg_tvalid && UG_rx_portg_tready && vacancy_cnt_q == 2'h1);
      la_rx_portf_tvalid_stg1_d = la_rx_portf_tvalid_stg1 &&
                                  !(LA_rx_portf_tvalid && UG_rx_portf_tready && vacancy_cnt_q == 2'h1);
      la_rx_porte_tvalid_stg1_d = la_rx_porte_tvalid_stg1 &&
                                  !(LA_rx_porte_tvalid && UG_rx_porte_tready && vacancy_cnt_q == 2'h1);
      la_rx_portd_tvalid_stg1_d = la_rx_portd_tvalid_stg1 &&
                                  !(LA_rx_portd_tvalid && UG_rx_portd_tready && vacancy_cnt_q == 2'h1);
      la_rx_portc_tvalid_stg1_d = la_rx_portc_tvalid_stg1 &&
                                  !(LA_rx_portc_tvalid && UG_rx_portc_tready && vacancy_cnt_q == 2'h1);
      la_rx_portb_tvalid_stg1_d = la_rx_portb_tvalid_stg1 &&
                                  !(LA_rx_portb_tvalid && UG_rx_portb_tready && vacancy_cnt_q == 2'h1);
      la_rx_porta_tvalid_stg1_d = la_rx_porta_tvalid_stg1 &&
                                  !(LA_rx_porta_tvalid && UG_rx_porta_tready && vacancy_cnt_q == 2'h1);

      // Stage 2 (contains both set and clear logic)
      la_rx_porth_tvalid_stg2_d = la_rx_porth_tvalid_stg2 &&
                                  !(LA_rx_porth_tvalid && UG_rx_porth_tready && vacancy_cnt_q == 2'h2);
      la_rx_portg_tvalid_stg2_d = la_rx_portg_tvalid_stg2 &&
                                  !(LA_rx_portg_tvalid && UG_rx_portg_tready && vacancy_cnt_q == 2'h2);
      la_rx_portf_tvalid_stg2_d = la_rx_portf_tvalid_stg2 &&
                                  !(LA_rx_portf_tvalid && UG_rx_portf_tready && vacancy_cnt_q == 2'h2);
      la_rx_porte_tvalid_stg2_d = la_rx_porte_tvalid_stg2 &&
                                  !(LA_rx_porte_tvalid && UG_rx_porte_tready && vacancy_cnt_q == 2'h2);
      la_rx_portd_tvalid_stg2_d = la_rx_portd_tvalid_stg2 &&
                                  !(LA_rx_portd_tvalid && UG_rx_portd_tready && vacancy_cnt_q == 2'h2);
      la_rx_portc_tvalid_stg2_d = la_rx_portc_tvalid_stg2 &&
                                  !(LA_rx_portc_tvalid && UG_rx_portc_tready && vacancy_cnt_q == 2'h2);
      la_rx_portb_tvalid_stg2_d = la_rx_portb_tvalid_stg2 &&
                                  !(LA_rx_portb_tvalid && UG_rx_portb_tready && vacancy_cnt_q == 2'h2);
      la_rx_porta_tvalid_stg2_d = la_rx_porta_tvalid_stg2 &&
                                  !(LA_rx_porta_tvalid && UG_rx_porta_tready && vacancy_cnt_q == 2'h2);
    end
  end
  // }}} End of Demux Logic ---------------


  // {{{ Port Interface Control -----------

  // final determination for TVALID
  assign la_rx_porta_tvalid_d = vacancy_cnt != 2'h0 && ~|(tvalid_list & 8'b01111111) &&
                                ((la_rx_porta_tvalid_stg0 && !la_rx_porta_any_tvalid_stg1) ||
                                 (la_rx_porta_tvalid_stg1 &&
                                   (vacancy_cnt_q == 2'h2 ||
                                   !(UG_rx_porta_tready && LA_rx_porta_tvalid && !la_rx_porta_any_tvalid_stg2))) ||
                                 (la_rx_porta_tvalid_stg2 && !(UG_rx_porta_tready && LA_rx_porta_tvalid)));
  assign la_rx_portb_tvalid_d = vacancy_cnt != 2'h0 && ~|(tvalid_list & 8'b10111111) &&
                                ((la_rx_portb_tvalid_stg0 && !la_rx_portb_any_tvalid_stg1) ||
                                 (la_rx_portb_tvalid_stg1 &&
                                   (vacancy_cnt_q == 2'h2 ||
                                   !(UG_rx_portb_tready && LA_rx_portb_tvalid && !la_rx_portb_any_tvalid_stg2))) ||
                                 (la_rx_portb_tvalid_stg2 && !(UG_rx_portb_tready && LA_rx_portb_tvalid)));
  assign la_rx_portc_tvalid_d = vacancy_cnt != 2'h0 && ~|(tvalid_list & 8'b11011111) &&
                                ((la_rx_portc_tvalid_stg0 && !la_rx_portc_any_tvalid_stg1) ||
                                 (la_rx_portc_tvalid_stg1 &&
                                   (vacancy_cnt_q == 2'h2 ||
                                   !(UG_rx_portc_tready && LA_rx_portc_tvalid && !la_rx_portc_any_tvalid_stg2))) ||
                                 (la_rx_portc_tvalid_stg2 && !(UG_rx_portc_tready && LA_rx_portc_tvalid)));
  assign la_rx_portd_tvalid_d = vacancy_cnt != 2'h0 && ~|(tvalid_list & 8'b11101111) &&
                                ((la_rx_portd_tvalid_stg0 && !la_rx_portd_any_tvalid_stg1) ||
                                 (la_rx_portd_tvalid_stg1 && 
                                   (vacancy_cnt_q == 2'h2 ||
                                   !(UG_rx_portd_tready && LA_rx_portd_tvalid && !la_rx_portd_any_tvalid_stg2))) ||
                                 (la_rx_portd_tvalid_stg2 && !(UG_rx_portd_tready && LA_rx_portd_tvalid)));
  assign la_rx_porte_tvalid_d = vacancy_cnt != 2'h0 && ~|(tvalid_list & 8'b11110111) &&
                                ((la_rx_porte_tvalid_stg0 && !la_rx_porte_any_tvalid_stg1) ||
                                 (la_rx_porte_tvalid_stg1 &&
                                   (vacancy_cnt_q == 2'h2 ||
                                   !(UG_rx_porte_tready && LA_rx_porte_tvalid && !la_rx_porte_any_tvalid_stg2))) ||
                                 (la_rx_porte_tvalid_stg2 && !(UG_rx_porte_tready && LA_rx_porte_tvalid)));
  assign la_rx_portf_tvalid_d = vacancy_cnt != 2'h0 && ~|(tvalid_list & 8'b11111011) &&
                                ((la_rx_portf_tvalid_stg0 && !la_rx_portf_any_tvalid_stg1) ||
                                 (la_rx_portf_tvalid_stg1 &&
                                   (vacancy_cnt_q == 2'h2 ||
                                   !(UG_rx_portf_tready && LA_rx_portf_tvalid && !la_rx_portf_any_tvalid_stg2))) ||
                                 (la_rx_portf_tvalid_stg2 && !(UG_rx_portf_tready && LA_rx_portf_tvalid)));
  assign la_rx_portg_tvalid_d = vacancy_cnt != 2'h0 && ~|(tvalid_list & 8'b11111101) &&
                                ((la_rx_portg_tvalid_stg0 && !la_rx_portg_any_tvalid_stg1) ||
                                 (la_rx_portg_tvalid_stg1 &&
                                   (vacancy_cnt_q == 2'h2 ||
                                   !(UG_rx_portg_tready && LA_rx_portg_tvalid && !la_rx_portg_any_tvalid_stg2))) ||
                                 (la_rx_portg_tvalid_stg2 && !(UG_rx_portg_tready && LA_rx_portg_tvalid)));
  assign la_rx_porth_tvalid_d = vacancy_cnt != 2'h0 && ~|(tvalid_list & 8'b11111110) &&
                                ((la_rx_porth_tvalid_stg0 && !la_rx_porth_any_tvalid_stg1) ||
                                 (la_rx_porth_tvalid_stg1 &&
                                   (vacancy_cnt_q == 2'h2 ||
                                   !(UG_rx_porth_tready && LA_rx_porth_tvalid && !la_rx_porth_any_tvalid_stg2))) ||
                                 (la_rx_porth_tvalid_stg2 && !(UG_rx_porth_tready && LA_rx_porth_tvalid)));


  // final determination for TLAST
  assign la_rx_porta_tlast_d =
          la_rx_porta_tvalid_stg2 && !(UG_rx_porta_tready && LA_rx_porta_tvalid) ? le_lhrx_tlast_stg2 :
          la_rx_porta_tvalid_stg2 && UG_rx_porta_tready && LA_rx_porta_tvalid    ? le_lhrx_tlast_stg1 :
          la_rx_porta_tvalid_stg1 && !(UG_rx_porta_tready && LA_rx_porta_tvalid) ? le_lhrx_tlast_stg1 :
          la_rx_porta_tvalid_stg1 && UG_rx_porta_tready && LA_rx_porta_tvalid    ? le_lhrx_tlast_q    :
          la_rx_porta_tvalid_stg0                                                ? le_lhrx_tlast_q    :  1'b0;
  assign la_rx_portb_tlast_d =
          la_rx_portb_tvalid_stg2 && !(UG_rx_portb_tready && LA_rx_portb_tvalid) ? le_lhrx_tlast_stg2 :
          la_rx_portb_tvalid_stg2 && UG_rx_portb_tready && LA_rx_portb_tvalid    ? le_lhrx_tlast_stg1 :
          la_rx_portb_tvalid_stg1 && !(UG_rx_portb_tready && LA_rx_portb_tvalid) ? le_lhrx_tlast_stg1 :
          la_rx_portb_tvalid_stg1 && UG_rx_portb_tready && LA_rx_portb_tvalid    ? le_lhrx_tlast_q    :
          la_rx_portb_tvalid_stg0                                                ? le_lhrx_tlast_q    :  1'b0;
  assign la_rx_portc_tlast_d =
          la_rx_portc_tvalid_stg2 && !(UG_rx_portc_tready && LA_rx_portc_tvalid) ? le_lhrx_tlast_stg2 :
          la_rx_portc_tvalid_stg2 && UG_rx_portc_tready && LA_rx_portc_tvalid    ? le_lhrx_tlast_stg1 :
          la_rx_portc_tvalid_stg1 && !(UG_rx_portc_tready && LA_rx_portc_tvalid) ? le_lhrx_tlast_stg1 :
          la_rx_portc_tvalid_stg1 && UG_rx_portc_tready && LA_rx_portc_tvalid    ? le_lhrx_tlast_q    :
          la_rx_portc_tvalid_stg0                                                ? le_lhrx_tlast_q    :  1'b0;
  assign la_rx_portd_tlast_d =
          la_rx_portd_tvalid_stg2 && !(UG_rx_portd_tready && LA_rx_portd_tvalid) ? le_lhrx_tlast_stg2 :
          la_rx_portd_tvalid_stg2 && UG_rx_portd_tready && LA_rx_portd_tvalid    ? le_lhrx_tlast_stg1 :
          la_rx_portd_tvalid_stg1 && !(UG_rx_portd_tready && LA_rx_portd_tvalid) ? le_lhrx_tlast_stg1 :
          la_rx_portd_tvalid_stg1 && UG_rx_portd_tready && LA_rx_portd_tvalid    ? le_lhrx_tlast_q    :
          la_rx_portd_tvalid_stg0                                                ? le_lhrx_tlast_q    :  1'b0;
  assign la_rx_porte_tlast_d =
          la_rx_porte_tvalid_stg2 && !(UG_rx_porte_tready && LA_rx_porte_tvalid) ? le_lhrx_tlast_stg2 :
          la_rx_porte_tvalid_stg2 && UG_rx_porte_tready && LA_rx_porte_tvalid    ? le_lhrx_tlast_stg1 :
          la_rx_porte_tvalid_stg1 && !(UG_rx_porte_tready && LA_rx_porte_tvalid) ? le_lhrx_tlast_stg1 :
          la_rx_porte_tvalid_stg1 && UG_rx_porte_tready && LA_rx_porte_tvalid    ? le_lhrx_tlast_q    :
          la_rx_porte_tvalid_stg0                                                ? le_lhrx_tlast_q    :  1'b0;
  assign la_rx_portf_tlast_d =
          la_rx_portf_tvalid_stg2 && !(UG_rx_portf_tready && LA_rx_portf_tvalid) ? le_lhrx_tlast_stg2 :
          la_rx_portf_tvalid_stg2 && UG_rx_portf_tready && LA_rx_portf_tvalid    ? le_lhrx_tlast_stg1 :
          la_rx_portf_tvalid_stg1 && !(UG_rx_portf_tready && LA_rx_portf_tvalid) ? le_lhrx_tlast_stg1 :
          la_rx_portf_tvalid_stg1 && UG_rx_portf_tready && LA_rx_portf_tvalid    ? le_lhrx_tlast_q    :
          la_rx_portf_tvalid_stg0                                                ? le_lhrx_tlast_q    :  1'b0;
  assign la_rx_portg_tlast_d =
          la_rx_portg_tvalid_stg2 && !(UG_rx_portg_tready && LA_rx_portg_tvalid) ? le_lhrx_tlast_stg2 :
          la_rx_portg_tvalid_stg2 && UG_rx_portg_tready && LA_rx_portg_tvalid    ? le_lhrx_tlast_stg1 :
          la_rx_portg_tvalid_stg1 && !(UG_rx_portg_tready && LA_rx_portg_tvalid) ? le_lhrx_tlast_stg1 :
          la_rx_portg_tvalid_stg1 && UG_rx_portg_tready && LA_rx_portg_tvalid    ? le_lhrx_tlast_q    :
          la_rx_portg_tvalid_stg0                                                ? le_lhrx_tlast_q    :  1'b0;
  assign la_rx_porth_tlast_d =
          la_rx_porth_tvalid_stg2 && !(UG_rx_porth_tready && LA_rx_porth_tvalid) ? le_lhrx_tlast_stg2 :
          la_rx_porth_tvalid_stg2 && UG_rx_porth_tready && LA_rx_porth_tvalid    ? le_lhrx_tlast_stg1 :
          la_rx_porth_tvalid_stg1 && !(UG_rx_porth_tready && LA_rx_porth_tvalid) ? le_lhrx_tlast_stg1 :
          la_rx_porth_tvalid_stg1 && UG_rx_porth_tready && LA_rx_porth_tvalid    ? le_lhrx_tlast_q    :
          la_rx_porth_tvalid_stg0                                                ? le_lhrx_tlast_q    :  1'b0;


  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LA_rx_porta_tvalid <= #TCQ 1'b0;
      LA_rx_portb_tvalid <= #TCQ 1'b0;
      LA_rx_portc_tvalid <= #TCQ 1'b0;
      LA_rx_portd_tvalid <= #TCQ 1'b0;
      LA_rx_porte_tvalid <= #TCQ 1'b0;
      LA_rx_portf_tvalid <= #TCQ 1'b0;
      LA_rx_portg_tvalid <= #TCQ 1'b0;
      LA_rx_porth_tvalid <= #TCQ 1'b0;

      LA_rx_porta_tlast  <= #TCQ 1'b0;
      LA_rx_portb_tlast  <= #TCQ 1'b0;
      LA_rx_portc_tlast  <= #TCQ 1'b0;
      LA_rx_portd_tlast  <= #TCQ 1'b0;
      LA_rx_porte_tlast  <= #TCQ 1'b0;
      LA_rx_portf_tlast  <= #TCQ 1'b0;
      LA_rx_portg_tlast  <= #TCQ 1'b0;
      LA_rx_porth_tlast  <= #TCQ 1'b0;
    end else begin
      LA_rx_porta_tvalid <= #TCQ la_rx_porta_tvalid_d;
      LA_rx_portb_tvalid <= #TCQ la_rx_portb_tvalid_d;
      LA_rx_portc_tvalid <= #TCQ la_rx_portc_tvalid_d;
      LA_rx_portd_tvalid <= #TCQ la_rx_portd_tvalid_d;
      LA_rx_porte_tvalid <= #TCQ la_rx_porte_tvalid_d;
      LA_rx_portf_tvalid <= #TCQ la_rx_portf_tvalid_d;
      LA_rx_portg_tvalid <= #TCQ la_rx_portg_tvalid_d;
      LA_rx_porth_tvalid <= #TCQ la_rx_porth_tvalid_d;

      LA_rx_porta_tlast  <= #TCQ la_rx_porta_tlast_d;
      LA_rx_portb_tlast  <= #TCQ la_rx_portb_tlast_d;
      LA_rx_portc_tlast  <= #TCQ la_rx_portc_tlast_d;
      LA_rx_portd_tlast  <= #TCQ la_rx_portd_tlast_d;
      LA_rx_porte_tlast  <= #TCQ la_rx_porte_tlast_d;
      LA_rx_portf_tlast  <= #TCQ la_rx_portf_tlast_d;
      LA_rx_portg_tlast  <= #TCQ la_rx_portg_tlast_d;
      LA_rx_porth_tlast  <= #TCQ la_rx_porth_tlast_d;
    end
  end

  // TREADY generation - if data is sitting on the port to the user and has
  // not been accepted, we cannot accept the next beat of data.
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      la_lhrx_tready_d <= #TCQ 1'b0;
    end else begin
      if (clear_on_error) begin
        la_lhrx_tready_d <= #TCQ !le_out_of_packet_lhrx_q;
      end else begin
        la_lhrx_tready_d <= #TCQ vacancy_cnt < 2'h2 || |(tready_list & tvalid_list);
      end
    end
  end


  assign vacancy_cnt = (lhrx_advance_unqual) + (la_rx_port_any_tvalid_stg1) +
                       (la_rx_port_any_tvalid_stg2) - |(tready_list & tvalid_list);

  // Error detection logic
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LA_port_decode_error <= #TCQ 1'b0;
      vacancy_cnt_q        <= #TCQ 2'h0;
      clear_on_error       <= #TCQ 1'b0;
    end else begin
      LA_port_decode_error <= #TCQ port_decode_error_d;
      vacancy_cnt_q  <= #TCQ vacancy_cnt;
      if (le_out_of_packet_lhrx_q) begin
        clear_on_error       <= #TCQ 1'b0;
      end else if (port_decode_error_d) begin
        clear_on_error       <= #TCQ 1'b1;
      end
    end
  end

  // }}} End of Port Interface Control ----


  // {{{ Coverage and Assertions ----------

    // *- COVERAGE (cp_LAR_parameter_configurations)
    // Observe an agreed-upon set of parameter configurations

    // *- COVERAGE (cp_LAR_port_1_hit)
    // Observe one and only one port get a hit on a packet

    // *- COVERAGE (cp_LAR_port_2_hit)
    // Observe two ports get a hit on the same packet

    // *- COVERAGE (cp_LAR_port_3_hit)
    // Observe three ports get a hit on the same packet

    // *- COVERAGE (cp_LAR_port_no_hit)
    // Observe a packet that hits none of the ports with FALL_THROUGH set and unset

    // *- ASSERTION (ap_LAR_tvalid_behavior)
    // Only one TVALID from the RX Arbiter may ever be asserted

    // *- COVERAGE (cp_LAR_tready_drop_first)
    // Observe a destination's TREADY drop on the first beat of a packet

    // *- COVERAGE (cp_LAR_tready_drop_last)
    // Observe a destination's TREADY drop on the last beat of a packet

    // *- COVERAGE (cp_LAR_tready_drop_mid)
    // Observe a destination's TREADY drop on the middle of a packet

    // *- COVERAGE (cp_LAR_back_to_back_same_dest)
    // Observe back-to-back packets going to the same destination

    // *- COVERAGE (cp_LAR_back_to_back_different_dest)
    // Observe back-to-back packets going to different destinations

    // *- COVERAGE (cp_LAR_back_to_back_different_dest_2)
    // Observe back-to-back packets going to different destinations,
    // where the second packet could have gone to the first destination
    // if not for stricter criteria

    // *- COVERAGE (cp_LAR_tvalid_drop_second)
    // Observe the header encoder drop its TVALID after the first valid beat

    // *- COVERAGE (cp_LAR_tvalid_drop_last)
    // Observe the header encoder drop its TVALID one cycle before the last beat

    // *- COVERAGE (cp_LAR_tvalid_drop_mid)
    // Observe the header encoder drop TVALID in the middle of a packet

    // *- COVERAGE (cp_LAR_all_hits)
    // Cover hits of every type: FTYPE[1:5], TTYPE[1:5], STAT[1:2], LCSBA

    // *- COVERAGE (cp_LAR_partial_hit)
    // Observe a partial match - FTYPE but not TTYPE, TTYPE but not FTYPE

    // *- COVERAGE (cp_LAR_portx_tvalid_d)
    // Observe a specific logic sequence for portx_tvalid_d that was added
    // for v1.4 as a result of a customer bug:
    // !(la_rx_port*_tvalid_stg0 && !la_rx_port*_any_tvalid_stg1) &&
    // (la_rx_port*_tvalid_stg1 && vacancy_cnt_q == 2'h2)

  // }}} End Coverage and Assertions -------------


endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/log/log_arb/srio_gen2_v4_1_16_arb_tx.v#3 $
//
//----------------------------------------------------------------------
//
// ARB_TX
// Description:
// This module holds the transmit logic for the Arbiter
//
// Hierarchy:
// LOG_TOP
//    |_____ARB_TX <-- this module
//             |_____ARB_TX_USER_IF
//             |_____ARB_TX_MUX
//             |_____EVAL_LOG_CLK
//    |_____ARB_RX
// ---------------------------------------------------------------------

`timescale 1ps/1ps

// ------------------------------------------------
// below attribute is added to supress the synthesis warnings in vivado tool 8:3332
(* DowngradeIPIdentifiedWarnings="yes" *)
// ------------------------------------------------

module srio_gen2_v4_1_16_arb_tx



  #(
   // {{{ Parameter declarations -----------
    parameter TCQ                     = 100,  // in pS
    parameter EVAL                    = 1,    // Includes the evaluation timer

    parameter TX_ENABLE_FAIRNESS      = 1,    // When set, use tiebreaking technique {0,1}

    parameter TX_PORTA_HELLO          = 1,    // When set, HELLO format is in use {0,1}
    parameter TX_PORTB_HELLO          = 1,    // When set, HELLO format is in use {0,1}
    parameter TX_PORTC_HELLO          = 1,    // When set, HELLO format is in use {0,1}
    parameter TX_PORTD_HELLO          = 1,    // When set, HELLO format is in use {0,1}
    parameter TX_PORTE_HELLO          = 1,    // When set, HELLO format is in use {0,1}
    parameter TX_PORTF_HELLO          = 1,    // When set, HELLO format is in use {0,1}
    parameter TX_PORTG_HELLO          = 1,    // When set, HELLO format is in use {0,1}
    parameter TX_PORTH_HELLO          = 1,    // When set, HELLO format is in use {0,1}

    parameter TX_PORTA_ENABLE         = 1,    // Indicates if a port is enabled {0,1}
    parameter TX_PORTB_ENABLE         = 1,    // Indicates if a port is enabled {0,1}
    parameter TX_PORTC_ENABLE         = 1,    // Indicates if a port is enabled {0,1}
    parameter TX_PORTD_ENABLE         = 1,    // Indicates if a port is enabled {0,1}
    parameter TX_PORTE_ENABLE         = 1,    // Indicates if a port is enabled {0,1}
    parameter TX_PORTF_ENABLE         = 1,    // Indicates if a port is enabled {0,1}
    parameter TX_PORTG_ENABLE         = 1,    // Indicates if a port is enabled {0,1}
    parameter TX_PORTH_ENABLE         = 1,    // Indicates if a port is enabled {0,1}

    parameter TX_PORTA_PRIORITY       = 1,    // Indicates the priority of a port {0-3}
    parameter TX_PORTB_PRIORITY       = 1,    // Indicates the priority of a port {0-3}
    parameter TX_PORTC_PRIORITY       = 1,    // Indicates the priority of a port {0-3}
    parameter TX_PORTD_PRIORITY       = 1,    // Indicates the priority of a port {0-3}
    parameter TX_PORTE_PRIORITY       = 1,    // Indicates the priority of a port {0-3}
    parameter TX_PORTF_PRIORITY       = 1,    // Indicates the priority of a port {0-3}
    parameter TX_PORTG_PRIORITY       = 1,    // Indicates the priority of a port {0-3}
    parameter TX_PORTH_PRIORITY       = 1,    // Indicates the priority of a port {0-3}

    parameter TX_PORTA_RESP_CLASS     = 0,    // When set, indicates a Response interface {0,1}
    parameter TX_PORTB_RESP_CLASS     = 0,    // When set, indicates a Response interface {0,1}
    parameter TX_PORTC_RESP_CLASS     = 0,    // When set, indicates a Response interface {0,1}
    parameter TX_PORTD_RESP_CLASS     = 0,    // When set, indicates a Response interface {0,1}
    parameter TX_PORTE_RESP_CLASS     = 0,    // When set, indicates a Response interface {0,1}
    parameter TX_PORTF_RESP_CLASS     = 0,    // When set, indicates a Response interface {0,1}
    parameter TX_PORTG_RESP_CLASS     = 0,    // When set, indicates a Response interface {0,1}
    parameter TX_PORTH_RESP_CLASS     = 0,    // When set, indicates a Response interface {0,1}
    parameter CRF_SUPPORT             = 1)      

   // }}} ----------------------------------
   (
   // {{{ port declarations ----------------
    // clocks and resets and general signals
    input             log_clk,                // PHY interface clock
    input             log_rst,                // Reset for PHY clock Domain

    // PORTA TX Interface
    input             UG_tx_porta_tvalid,     // Valid Packet Beat
    output            LA_tx_porta_tready,     // Packet Beat Accepted
    input      [63:0] UG_tx_porta_tdata,      // Packet Data
    input       [7:0] UG_tx_porta_tkeep,      // Valid bytes in this beat, only valid on last
    input             UG_tx_porta_tlast,      // Last Beat
    input      [39:0] UG_tx_porta_tuser,      // {DEST_ID, SRC_ID, 5'h0, VC, CRF, 1'b0}

    // PORTB TX Interface
    input             UG_tx_portb_tvalid,     // Valid Packet Beat
    output            LA_tx_portb_tready,     // Packet Beat Accepted
    input      [63:0] UG_tx_portb_tdata,      // Packet Data
    input       [7:0] UG_tx_portb_tkeep,      // Valid bytes in this beat, only valid on last
    input             UG_tx_portb_tlast,      // Last Beat
    input      [39:0] UG_tx_portb_tuser,      // {DEST_ID, SRC_ID, 5'h0, VC, CRF, 1'b0}

    // PORTC TX Interface
    input             UG_tx_portc_tvalid,     // Valid Packet Beat
    output            LA_tx_portc_tready,     // Packet Beat Accepted
    input      [63:0] UG_tx_portc_tdata,      // Packet Data
    input       [7:0] UG_tx_portc_tkeep,      // Valid bytes in this beat, only valid on last
    input             UG_tx_portc_tlast,      // Last Beat
    input      [39:0] UG_tx_portc_tuser,      // {DEST_ID, SRC_ID, 5'h0, VC, CRF, 1'b0}

    // PORTD TX Interface
    input             UG_tx_portd_tvalid,     // Valid Packet Beat
    output            LA_tx_portd_tready,     // Packet Beat Accepted
    input      [63:0] UG_tx_portd_tdata,      // Packet Data
    input       [7:0] UG_tx_portd_tkeep,      // Valid bytes in this beat, only valid on last
    input             UG_tx_portd_tlast,      // Last Beat
    input      [39:0] UG_tx_portd_tuser,      // {DEST_ID, SRC_ID, 5'h0, VC, CRF, 1'b0}

    // PORTE TX Interface
    input             UG_tx_porte_tvalid,     // Valid Packet Beat
    output            LA_tx_porte_tready,     // Packet Beat Accepted
    input      [63:0] UG_tx_porte_tdata,      // Packet Data
    input       [7:0] UG_tx_porte_tkeep,      // Valid bytes in this beat, only valid on last
    input             UG_tx_porte_tlast,      // Last Beat
    input      [39:0] UG_tx_porte_tuser,      // {DEST_ID, SRC_ID, 5'h0, VC, CRF, 1'b0}

    // PORTF TX Interface
    input             UG_tx_portf_tvalid,     // Valid Packet Beat
    output            LA_tx_portf_tready,     // Packet Beat Accepted
    input      [63:0] UG_tx_portf_tdata,      // Packet Data
    input       [7:0] UG_tx_portf_tkeep,      // Valid bytes in this beat, only valid on last
    input             UG_tx_portf_tlast,      // Last Beat
    input      [39:0] UG_tx_portf_tuser,      // {DEST_ID, SRC_ID, 5'h0, VC, CRF, 1'b0}

    // PORTG TX Interface
    input             UG_tx_portg_tvalid,     // Valid Packet Beat
    output            LA_tx_portg_tready,     // Packet Beat Accepted
    input      [63:0] UG_tx_portg_tdata,      // Packet Data
    input       [7:0] UG_tx_portg_tkeep,      // Valid bytes in this beat, only valid on last
    input             UG_tx_portg_tlast,      // Last Beat
    input      [39:0] UG_tx_portg_tuser,      // {DEST_ID, SRC_ID, 5'h0, VC, CRF, 1'b0}

    // PORTH TX Interface
    input             UG_tx_porth_tvalid,     // Valid Packet Beat
    output            LA_tx_porth_tready,     // Packet Beat Accepted
    input      [63:0] UG_tx_porth_tdata,      // Packet Data
    input       [7:0] UG_tx_porth_tkeep,      // Valid bytes in this beat, only valid on last
    input             UG_tx_porth_tlast,      // Last Beat
    input      [39:0] UG_tx_porth_tuser,      // {DEST_ID, SRC_ID, 5'h0, VC, CRF, 1'b0}


    // Header Encoder TX Interface
    output            LA_lhtx_tvalid,         // Valid Packet Beat
    input             LD_lhtx_tready,         // Packet Beat Accepted
    output     [63:0] LA_lhtx_tdata,          // Packet Data
    output      [7:0] LA_lhtx_tkeep,          // Valid bytes in this beat, only valid on last
    output            LA_lhtx_tlast,          // Last Beat
    output     [39:0] LA_lhtx_tuser,          // {DEST_ID, SRC_ID, 3'h0, RESPONSE, HELLO_FMT, VC, CRF, 1'b0}

    // TX Buffer Interface
    input             BT_response_only,       // Buffer only has room for Resp Packets

    // Configuration signals
    input             PC_maint_only           // LOG can only send maint transactions

   // }}} ----------------------------------
   );


  // {{{ local parameters -----------------

  // Bit widths of each interface bus
  localparam PORT_ID      = 4;
  localparam TDATA_WIDTH  = 64;
  localparam TKEEP_WIDTH  = 8;
  localparam TUSER_WIDTH  = 40;
  localparam HELLO_BIT    = 1;
  localparam TREADY_WIDTH = 1;
  localparam TLAST_WIDTH  = 1;
  localparam TVALID_WIDTH = 1;
  localparam RESP_BIT     = 1; // currently not used

  // most of the data ports coming from interfaces are just considered data.
  // Add them to a large object for easier transport
  localparam TX_OBJECT_WIDTH = PORT_ID + TDATA_WIDTH + TKEEP_WIDTH + TUSER_WIDTH +
                               HELLO_BIT + TREADY_WIDTH + TLAST_WIDTH + TVALID_WIDTH;

  // move the parameters into an array, to be managed by a generate-for loop
  // parameters can't be two-dimensional. make it flat and bit-select later
  localparam [7:0] TX_PORT_HELLO = {TX_PORTH_HELLO[0], TX_PORTG_HELLO[0], TX_PORTF_HELLO[0],
                                    TX_PORTE_HELLO[0], TX_PORTD_HELLO[0], TX_PORTC_HELLO[0],
                                    TX_PORTB_HELLO[0], TX_PORTA_HELLO[0]}; 

  localparam [7:0] TX_PORT_RESP_CLASS = {TX_PORTH_RESP_CLASS[0], TX_PORTG_RESP_CLASS[0], TX_PORTF_RESP_CLASS[0],
                                         TX_PORTE_RESP_CLASS[0], TX_PORTD_RESP_CLASS[0], TX_PORTC_RESP_CLASS[0],
                                         TX_PORTB_RESP_CLASS[0], TX_PORTA_RESP_CLASS[0]};


  // count how many ports are going to each priority-based arbiter
  localparam [7:0] PRIO0_DEPTH = (TX_PORTA_ENABLE && TX_PORTA_PRIORITY == 0) +
                                 (TX_PORTB_ENABLE && TX_PORTB_PRIORITY == 0) +
                                 (TX_PORTC_ENABLE && TX_PORTC_PRIORITY == 0) +
                                 (TX_PORTD_ENABLE && TX_PORTD_PRIORITY == 0) +
                                 (TX_PORTE_ENABLE && TX_PORTE_PRIORITY == 0) +
                                 (TX_PORTF_ENABLE && TX_PORTF_PRIORITY == 0) +
                                 (TX_PORTG_ENABLE && TX_PORTG_PRIORITY == 0) +
                                 (TX_PORTH_ENABLE && TX_PORTH_PRIORITY == 0);

  localparam [7:0] PRIO1_DEPTH = (TX_PORTA_ENABLE && TX_PORTA_PRIORITY == 1) +
                                 (TX_PORTB_ENABLE && TX_PORTB_PRIORITY == 1) +
                                 (TX_PORTC_ENABLE && TX_PORTC_PRIORITY == 1) +
                                 (TX_PORTD_ENABLE && TX_PORTD_PRIORITY == 1) +
                                 (TX_PORTE_ENABLE && TX_PORTE_PRIORITY == 1) +
                                 (TX_PORTF_ENABLE && TX_PORTF_PRIORITY == 1) +
                                 (TX_PORTG_ENABLE && TX_PORTG_PRIORITY == 1) +
                                 (TX_PORTH_ENABLE && TX_PORTH_PRIORITY == 1);
  
  localparam [7:0] PRIO2_DEPTH = (TX_PORTA_ENABLE && TX_PORTA_PRIORITY == 2) +
                                 (TX_PORTB_ENABLE && TX_PORTB_PRIORITY == 2) +
                                 (TX_PORTC_ENABLE && TX_PORTC_PRIORITY == 2) +
                                 (TX_PORTD_ENABLE && TX_PORTD_PRIORITY == 2) +
                                 (TX_PORTE_ENABLE && TX_PORTE_PRIORITY == 2) +
                                 (TX_PORTF_ENABLE && TX_PORTF_PRIORITY == 2) +
                                 (TX_PORTG_ENABLE && TX_PORTG_PRIORITY == 2) +
                                 (TX_PORTH_ENABLE && TX_PORTH_PRIORITY == 2);
  
  localparam [7:0] PRIO3_DEPTH = (TX_PORTA_ENABLE && TX_PORTA_PRIORITY == 3) +
                                 (TX_PORTB_ENABLE && TX_PORTB_PRIORITY == 3) +
                                 (TX_PORTC_ENABLE && TX_PORTC_PRIORITY == 3) +
                                 (TX_PORTD_ENABLE && TX_PORTD_PRIORITY == 3) +
                                 (TX_PORTE_ENABLE && TX_PORTE_PRIORITY == 3) +
                                 (TX_PORTF_ENABLE && TX_PORTF_PRIORITY == 3) +
                                 (TX_PORTG_ENABLE && TX_PORTG_PRIORITY == 3) +
                                 (TX_PORTH_ENABLE && TX_PORTH_PRIORITY == 3);

  // put the values into a bus to use in the generate-for loop
  // params can't be two-dimensional, must use bit select later
  localparam [31:0] PRIO_DEPTH = {PRIO3_DEPTH, PRIO2_DEPTH, PRIO1_DEPTH, PRIO0_DEPTH};

  // dedicated maintenance ports are G and H.
  // If more flexibility is required, make into a param
  localparam [7:0] MAINT_PORTS = {1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};

  // unique identifiers for each physical port
  localparam PORTA = 4'h0;
  localparam PORTB = 4'h1;
  localparam PORTC = 4'h2;
  localparam PORTD = 4'h3;
  localparam PORTE = 4'h4;
  localparam PORTF = 4'h5;
  localparam PORTG = 4'h6;
  localparam PORTH = 4'h7;
  localparam NONE  = 4'hF;

  // }}} End local parameters -------------


  // {{{ wire declarations ----------------

  // pre pipeline results
  wire [63:0]  la_lhtx_tdata_pre;
  wire  [7:0]  la_lhtx_tkeep_pre;
  wire [39:0]  la_lhtx_tuser_pre;
  wire         la_lhtx_tlast_pre;
  wire         la_lhtx_tvalid_pre;
  wire         ld_lhtx_tready_pre;

  // common-use signals
  reg         log_rst_q = 1;           // Registered reset signal
  reg         log_packet_first_beat;   // * This is the eval timeout signal *
  wire        log_packet_first_beat_d; // * This is the eval timeout signal *
  reg         bt_response_only_q;      // registered version of respose-only signal
  reg         pc_maint_only_q;         // registered version of maint-only signal
  wire [7:0]  port_tvalid_mod;         // qualify the valid signal from the user to ignore the user in certain cases
  reg  [7:0]  port_tvalid_mod_q;       // Registered port_tvalid_mod
  wire [7:0]  la_port_mask_tvalid;     // when set, enables tvalid to propigate
  reg  [7:0]  disable_packet;
  reg  [7:0]  disable_packet_q;


  // result of the registered user interface
  // put into arrays for easier transport and use in generates
  // simple assignment - [0] is porta, [1] is portb, etc.
  reg   [7:0] la_tx_port_tready_d;
  reg   [7:0] la_tx_port_tready_dd;
  wire  [7:0] ug_tx_port_tvalid_q;
  wire  [7:0] ug_tx_port_tvalid_raw_q;
  wire [63:0] ug_tx_port_tdata_q  [7:0];
  wire  [7:0] ug_tx_port_tkeep_q  [7:0];
  wire  [7:0] ug_tx_port_tlast_q;
  wire [39:0] ug_tx_port_tuser_q  [7:0];

  wire  [7:0] la_tx_port_tready;
  wire  [7:0] ug_tx_port_tvalid;
  wire [63:0] ug_tx_port_tdata  [7:0];
  wire  [7:0] ug_tx_port_tkeep  [7:0];
  wire  [7:0] ug_tx_port_tlast;
  wire [39:0] ug_tx_port_tuser  [7:0];

  wire        la_no_advance     = la_lhtx_tvalid_pre && !ld_lhtx_tready_pre;
  wire        advance_condition = ld_lhtx_tready_pre || !la_lhtx_tvalid_pre;

  // create object blocks for simplicity of transfer. Each physical port has an associated object
  wire [TX_OBJECT_WIDTH-1:0] port_object_in [7:0];
  wire  [7:0]                port_object_last_beat;


  reg  [TX_OBJECT_WIDTH-1:0] winning_port_object;
  reg  [TX_OBJECT_WIDTH-1:0] winning_port_object_d;
  wire [TX_OBJECT_WIDTH-1:0] winning_port_object_dd;


  // individual priority winners and final winner
  wire [3:0]         port_winner_bus [PORT_ID-1:0];
  wire [PORT_ID-1:0] p0_port_winner = port_winner_bus[0];
  wire [PORT_ID-1:0] p1_port_winner = port_winner_bus[1];
  wire [PORT_ID-1:0] p2_port_winner = port_winner_bus[2];
  wire [PORT_ID-1:0] p3_port_winner = port_winner_bus[3];
  reg  [PORT_ID-1:0] port_winner;

  // TREADY combinatorial indicators
  reg la_tx_porta_tready_early;
  reg la_tx_portb_tready_early;
  reg la_tx_portc_tready_early;
  reg la_tx_portd_tready_early;
  reg la_tx_porte_tready_early;
  reg la_tx_portf_tready_early;
  reg la_tx_portg_tready_early;
  reg la_tx_porth_tready_early;

  // }}} End wire declarations ------------


  // {{{ Reset Structure ------------------

  // by rule, we must register the resets before we use them. This is not a
  // synchronizing circuit but rather a method to reduce fanout on the resets.
  always @(posedge log_clk or posedge log_rst) begin
    if (log_rst)
      log_rst_q <= #TCQ 1'b1;
    else
      log_rst_q <= #TCQ 1'b0;
  end

  // }}} End of Reset Structure -----------


  // {{{ User Interface Registering -------

  // register each port interface
  //____________________________________________________________________________
  assign LA_tx_porta_tready   = la_tx_port_tready[0];
  assign ug_tx_port_tvalid[0] = UG_tx_porta_tvalid;
  assign ug_tx_port_tdata[0]  = UG_tx_porta_tdata;
  assign ug_tx_port_tkeep[0]  = UG_tx_porta_tkeep;
  assign ug_tx_port_tlast[0]  = UG_tx_porta_tlast;
  
  generate if (CRF_SUPPORT == 1) begin: porta_tuser_crf_en_gen
  assign ug_tx_port_tuser[0]  = UG_tx_porta_tuser;
  end endgenerate
  generate if (CRF_SUPPORT == 0) begin: porta_tuser_crf_dis_gen
       assign ug_tx_port_tuser[0]  = {UG_tx_porta_tuser[39:2],2'b0};
  end endgenerate
  //____________________________________________________________________________

  //____________________________________________________________________________
  assign LA_tx_portb_tready   = la_tx_port_tready[1];
  assign ug_tx_port_tvalid[1] = UG_tx_portb_tvalid;
  assign ug_tx_port_tdata[1]  = UG_tx_portb_tdata;
  assign ug_tx_port_tkeep[1]  = UG_tx_portb_tkeep;
  assign ug_tx_port_tlast[1]  = UG_tx_portb_tlast;
  generate if (CRF_SUPPORT == 1) begin: portb_tuser_crf_en_gen
  assign ug_tx_port_tuser[1]  = UG_tx_portb_tuser;
  end endgenerate
  generate if (CRF_SUPPORT == 0) begin: portb_tuser_crf_dis_gen
       assign ug_tx_port_tuser[1]  = {UG_tx_portb_tuser[39:2],2'b0};
  end endgenerate
  //____________________________________________________________________________

  //____________________________________________________________________________
  assign LA_tx_portc_tready   = la_tx_port_tready[2];
  assign ug_tx_port_tvalid[2] = UG_tx_portc_tvalid;
  assign ug_tx_port_tdata[2]  = UG_tx_portc_tdata;
  assign ug_tx_port_tkeep[2]  = UG_tx_portc_tkeep;
  assign ug_tx_port_tlast[2]  = UG_tx_portc_tlast;
  generate if (CRF_SUPPORT == 1) begin: portc_tuser_crf_en_gen
  assign ug_tx_port_tuser[2]  = UG_tx_portc_tuser;
  end endgenerate
  generate if (CRF_SUPPORT == 0) begin: portc_tuser_crf_dis_gen
       assign ug_tx_port_tuser[2]  = {UG_tx_portc_tuser[39:2],2'b0};
  end endgenerate
  //____________________________________________________________________________

  //____________________________________________________________________________
  assign LA_tx_portd_tready   = la_tx_port_tready[3];
  assign ug_tx_port_tvalid[3] = UG_tx_portd_tvalid;
  assign ug_tx_port_tdata[3]  = UG_tx_portd_tdata;
  assign ug_tx_port_tkeep[3]  = UG_tx_portd_tkeep;
  assign ug_tx_port_tlast[3]  = UG_tx_portd_tlast;
  generate if (CRF_SUPPORT == 1) begin: portd_tuser_crf_en_gen
  assign ug_tx_port_tuser[3]  = UG_tx_portd_tuser;
  end endgenerate
  generate if (CRF_SUPPORT == 0) begin: portd_tuser_crf_dis_gen
       assign ug_tx_port_tuser[3]  = {UG_tx_portd_tuser[39:2],2'b0};
  end endgenerate
  //____________________________________________________________________________

  //____________________________________________________________________________
  assign LA_tx_porte_tready   = la_tx_port_tready[4];
  assign ug_tx_port_tvalid[4] = UG_tx_porte_tvalid;
  assign ug_tx_port_tdata[4]  = UG_tx_porte_tdata;
  assign ug_tx_port_tkeep[4]  = UG_tx_porte_tkeep;
  assign ug_tx_port_tlast[4]  = UG_tx_porte_tlast;
  generate if (CRF_SUPPORT == 1) begin: porte_tuser_crf_en_gen
  assign ug_tx_port_tuser[4]  = UG_tx_porte_tuser;
  end endgenerate
  generate if (CRF_SUPPORT == 0) begin: porte_tuser_crf_dis_gen
       assign ug_tx_port_tuser[4]  = {UG_tx_porte_tuser[39:2],2'b0};
  end endgenerate
  //____________________________________________________________________________

  //____________________________________________________________________________
  assign LA_tx_portf_tready   = la_tx_port_tready[5];
  assign ug_tx_port_tvalid[5] = UG_tx_portf_tvalid;
  assign ug_tx_port_tdata[5]  = UG_tx_portf_tdata;
  assign ug_tx_port_tkeep[5]  = UG_tx_portf_tkeep;
  assign ug_tx_port_tlast[5]  = UG_tx_portf_tlast;
  generate if (CRF_SUPPORT == 1) begin: portf_tuser_crf_en_gen
  assign ug_tx_port_tuser[5]  = UG_tx_portf_tuser;
  end endgenerate
  generate if (CRF_SUPPORT == 0) begin: portf_tuser_crf_dis_gen
       assign ug_tx_port_tuser[5]  = {UG_tx_portf_tuser[39:2],2'b0};
  end endgenerate
  //____________________________________________________________________________

  //____________________________________________________________________________
  assign LA_tx_portg_tready   = la_tx_port_tready[6];
  assign ug_tx_port_tvalid[6] = UG_tx_portg_tvalid;
  assign ug_tx_port_tdata[6]  = UG_tx_portg_tdata;
  assign ug_tx_port_tkeep[6]  = UG_tx_portg_tkeep;
  assign ug_tx_port_tlast[6]  = UG_tx_portg_tlast;
  generate if (CRF_SUPPORT == 1) begin: portg_tuser_crf_en_gen
  assign ug_tx_port_tuser[6]  = UG_tx_portg_tuser;
  end endgenerate
  generate if (CRF_SUPPORT == 0) begin: portg_tuser_crf_dis_gen
       assign ug_tx_port_tuser[6]  = {UG_tx_portg_tuser[39:2],2'b0};
  end endgenerate
  //____________________________________________________________________________

  //____________________________________________________________________________
  assign LA_tx_porth_tready   = la_tx_port_tready[7];
  assign ug_tx_port_tvalid[7] = UG_tx_porth_tvalid;
  assign ug_tx_port_tdata[7]  = UG_tx_porth_tdata;
  assign ug_tx_port_tkeep[7]  = UG_tx_porth_tkeep;
  assign ug_tx_port_tlast[7]  = UG_tx_porth_tlast;
  generate if (CRF_SUPPORT == 1) begin: porth_tuser_crf_en_gen
  assign ug_tx_port_tuser[7]  = UG_tx_porth_tuser;
  end endgenerate
  generate if (CRF_SUPPORT == 0) begin: porth_tuser_crf_dis_gen
       assign ug_tx_port_tuser[7]  = {UG_tx_porth_tuser[39:2],2'b0};
  end endgenerate
  //____________________________________________________________________________

  // register the response_only signal, register the valid_mod signals
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      bt_response_only_q <= #TCQ 1'b0;
      pc_maint_only_q    <= #TCQ 1'b0;
      port_tvalid_mod_q  <= #TCQ 1'b0;
    end else begin
      bt_response_only_q <= #TCQ BT_response_only;
      pc_maint_only_q    <= #TCQ PC_maint_only;
      port_tvalid_mod_q  <= #TCQ ~disable_packet | (port_tvalid_mod & la_tx_port_tready_dd & 
                            {8{(!bt_response_only_q && BT_response_only) || (!pc_maint_only_q && PC_maint_only)}});
    end
  end
  assign la_port_mask_tvalid = ~disable_packet | (port_tvalid_mod & la_tx_port_tready_dd & 
                               {8{(!bt_response_only_q && BT_response_only) || (!pc_maint_only_q && PC_maint_only)}});


  // for loop used to instantiate the register ring between the user and core logic
  genvar jj;
  generate for (jj = 0; jj < 8; jj = jj+1) begin: user_if_gen
  reg out_of_packet, out_of_packet_q;

    srio_gen2_v4_1_16_arb_tx_user_if
      #(.TCQ                     (TCQ))
      arb_tx_user_if_port_inst
       (
        .log_clk                 (log_clk),
        .log_rst_q               (log_rst_q),

        .UG_tx_port_tvalid       (ug_tx_port_tvalid[jj]),
        .LA_tx_port_tready       (la_tx_port_tready[jj]),
        .UG_tx_port_tdata        (ug_tx_port_tdata[jj]),
        .UG_tx_port_tkeep        (ug_tx_port_tkeep[jj]),
        .UG_tx_port_tlast        (ug_tx_port_tlast[jj]),
        .UG_tx_port_tuser        (ug_tx_port_tuser[jj]),

        .LA_no_advance           (la_no_advance),
        .LA_port_mask_tvalid     (la_port_mask_tvalid[jj]),

        .UG_tx_port_tvalid_q     (ug_tx_port_tvalid_q[jj]),
        .UG_tx_port_tvalid_raw_q (ug_tx_port_tvalid_raw_q[jj]),
        .LA_tx_port_tready_d     (la_tx_port_tready_d[jj]),
        .UG_tx_port_tdata_q      (ug_tx_port_tdata_q[jj]),
        .UG_tx_port_tkeep_q      (ug_tx_port_tkeep_q[jj]),
        .UG_tx_port_tlast_q      (ug_tx_port_tlast_q[jj]),
        .UG_tx_port_tuser_q      (ug_tx_port_tuser_q[jj])
       );
  always @* begin
    out_of_packet           = out_of_packet_q    ;
    disable_packet[jj]      = disable_packet_q[jj];
    if (ug_tx_port_tlast_q[jj] && ug_tx_port_tvalid_raw_q[jj] && la_tx_port_tready_d[jj] && !la_no_advance) begin
      out_of_packet           = 1'b1;
      disable_packet[jj]      = (!TX_PORT_RESP_CLASS[jj] && BT_response_only) || (!MAINT_PORTS[jj] && PC_maint_only);
    end else if (port_tvalid_mod[jj] && la_tx_port_tready_d[jj]) begin
      out_of_packet           = 1'b0;
      disable_packet[jj]      = 1'b0;
    end else if (out_of_packet_q) begin
      disable_packet[jj]      = (!TX_PORT_RESP_CLASS[jj] && BT_response_only) || (!MAINT_PORTS[jj] && PC_maint_only);
    end
  end
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      out_of_packet_q       <= #TCQ 1'b1;
      disable_packet_q[jj]  <= #TCQ 1'b0;
    end else begin
      out_of_packet_q       <= #TCQ out_of_packet;
      disable_packet_q[jj]  <= #TCQ disable_packet[jj];
    end
  end

  assign port_tvalid_mod[jj] = ug_tx_port_tvalid_q[jj]; // && port_tvalid_mod_q[jj];
                               // resp/maint_only just asserted and the arbiter has already picked a winner
                               //((port_tvalid_mod_q[jj] && la_tx_port_tready_d[jj] && bt_rsp_maint_only_rose) ||
                               //(port_tvalid_mod_q[jj] || !disable_packet);

  assign port_object_in[jj] =
                             {jj, ug_tx_port_tdata_q[jj], ug_tx_port_tkeep_q[jj], ug_tx_port_tuser_q[jj],
                              TX_PORT_HELLO[jj] == 1, la_tx_port_tready_d[jj],
                              ug_tx_port_tlast_q[jj], port_tvalid_mod[jj]};
  assign port_object_last_beat[jj] = la_tx_port_tready_d[jj] && ug_tx_port_tlast_q[jj] && port_tvalid_mod[jj];

  end // for generate
  endgenerate

  // }}} End of User Interface Registering -


  // {{{ Priority 0 thru 3 Arbitration -----------
  // the for loop unrolls 4 time, one for each priority (0-3).
  genvar ii;
  generate for (ii = 0; ii < 4; ii = ii+1) begin: priority_arbitration_gen

    // Check to see if the number of ports for a given prio (PRIO_DEPTH) is non-zero
    if (PRIO_DEPTH[ii*8+:8] != 0) begin : prio_tx_arbiter

      reg  [TX_OBJECT_WIDTH-1:0] port1_object = 0;
      reg  [TX_OBJECT_WIDTH-1:0] port2_object = 0;
      reg  [TX_OBJECT_WIDTH-1:0] port3_object = 0;
      reg  [TX_OBJECT_WIDTH-1:0] port4_object = 0;
      reg  [TX_OBJECT_WIDTH-1:0] port5_object = 0;
      reg  [TX_OBJECT_WIDTH-1:0] port6_object = 0;
      reg  [TX_OBJECT_WIDTH-1:0] port7_object = 0;
      reg  [TX_OBJECT_WIDTH-1:0] port8_object = 0;

      // when these signals are set, it means that the interface port has been
      // assigned to an arbiter location already
      reg  portb_assigned;
      reg  portc_assigned;
      reg  portd_assigned;
      reg  porte_assigned;
      reg  portf_assigned;
      reg  portg_assigned;


      // this whole always block will be resolved before synthesis and costs nothing
      // in terms of resources. This procedure simply assigns ports to the appropriate
      // priority-based arbiter. Each port gets assigned in order from first to eighth (or last),
      // starting with port a and going to port h.
      always @* begin

        portb_assigned = 0;
        portc_assigned = 0;
        portd_assigned = 0;
        porte_assigned = 0;
        portf_assigned = 0;
        portg_assigned = 0;

        // first port assignment
        if (TX_PORTA_ENABLE && TX_PORTA_PRIORITY == ii) begin
          port1_object   = port_object_in[0];
        end else if (TX_PORTB_ENABLE && TX_PORTB_PRIORITY == ii) begin
          port1_object   = port_object_in[1];
          portb_assigned = 1;
        end else if (TX_PORTC_ENABLE && TX_PORTC_PRIORITY == ii) begin
          port1_object   = port_object_in[2];
          portc_assigned = 1;
        end else if (TX_PORTD_ENABLE && TX_PORTD_PRIORITY == ii) begin
          port1_object   = port_object_in[3];
          portd_assigned = 1;
        end else if (TX_PORTE_ENABLE && TX_PORTE_PRIORITY == ii) begin
          port1_object   = port_object_in[4];
          porte_assigned = 1;
        end else if (TX_PORTF_ENABLE && TX_PORTF_PRIORITY == ii) begin
          port1_object   = port_object_in[5];
          portf_assigned = 1;
        end else if (TX_PORTG_ENABLE && TX_PORTG_PRIORITY == ii) begin
          port1_object   = port_object_in[6];
          portg_assigned = 1;
        end else if (TX_PORTH_ENABLE && TX_PORTH_PRIORITY == ii) begin
          port1_object   = port_object_in[7];
        end else begin
          port1_object   = 'hx;
        end


        // second port assignment
        if (PRIO_DEPTH[ii*8+:8] > 1 && TX_PORTB_ENABLE && TX_PORTB_PRIORITY == ii && !portb_assigned) begin
          port2_object   = port_object_in[1];
        end else if (PRIO_DEPTH[ii*8+:8] > 1 && TX_PORTC_ENABLE && TX_PORTC_PRIORITY == ii && !portc_assigned) begin
          port2_object   = port_object_in[2];
          portc_assigned = 1;
        end else if (PRIO_DEPTH[ii*8+:8] > 1 && TX_PORTD_ENABLE && TX_PORTD_PRIORITY == ii && !portd_assigned) begin
          port2_object   = port_object_in[3];
          portd_assigned = 1;
        end else if (PRIO_DEPTH[ii*8+:8] > 1 && TX_PORTE_ENABLE && TX_PORTE_PRIORITY == ii && !porte_assigned) begin
          port2_object   = port_object_in[4];
          porte_assigned = 1;
        end else if (PRIO_DEPTH[ii*8+:8] > 1 && TX_PORTF_ENABLE && TX_PORTF_PRIORITY == ii && !portf_assigned) begin
          port2_object   = port_object_in[5];
          portf_assigned = 1;
        end else if (PRIO_DEPTH[ii*8+:8] > 1 && TX_PORTG_ENABLE && TX_PORTG_PRIORITY == ii && !portg_assigned) begin
          port2_object   = port_object_in[6];
          portg_assigned = 1;
        end else if (PRIO_DEPTH[ii*8+:8] > 1 && TX_PORTH_ENABLE && TX_PORTH_PRIORITY == ii) begin
          port2_object   = port_object_in[7];
        end else begin
          port2_object   = 'hx;
        end


        // third port assignment
        if (PRIO_DEPTH[ii*8+:8] > 2 && TX_PORTC_ENABLE && TX_PORTC_PRIORITY == ii && !portc_assigned) begin
          port3_object   = port_object_in[2];
        end else if (PRIO_DEPTH[ii*8+:8] > 2 && TX_PORTD_ENABLE && TX_PORTD_PRIORITY == ii && !portd_assigned) begin
          port3_object   = port_object_in[3];
          portd_assigned = 1;
        end else if (PRIO_DEPTH[ii*8+:8] > 2 && TX_PORTE_ENABLE && TX_PORTE_PRIORITY == ii && !porte_assigned) begin
          port3_object   = port_object_in[4];
          porte_assigned = 1;
        end else if (PRIO_DEPTH[ii*8+:8] > 2 && TX_PORTF_ENABLE && TX_PORTF_PRIORITY == ii && !portf_assigned) begin
          port3_object   = port_object_in[5];
          portf_assigned = 1;
        end else if (PRIO_DEPTH[ii*8+:8] > 2 && TX_PORTG_ENABLE && TX_PORTG_PRIORITY == ii && !portg_assigned) begin
          port3_object   = port_object_in[6];
          portg_assigned = 1;
        end else if (PRIO_DEPTH[ii*8+:8] > 2 && TX_PORTH_ENABLE && TX_PORTH_PRIORITY == ii) begin
          port3_object   = port_object_in[7];
        end else begin
          port3_object   = 'hx;
        end


        // fourth port assignment
        if (PRIO_DEPTH[ii*8+:8] > 3 && TX_PORTD_ENABLE && TX_PORTD_PRIORITY == ii && !portd_assigned) begin
          port4_object   = port_object_in[3];
        end else if (PRIO_DEPTH[ii*8+:8] > 3 && TX_PORTE_ENABLE && TX_PORTE_PRIORITY == ii && !porte_assigned) begin
          port4_object   = port_object_in[4];
          porte_assigned = 1;
        end else if (PRIO_DEPTH[ii*8+:8] > 3 && TX_PORTF_ENABLE && TX_PORTF_PRIORITY == ii && !portf_assigned) begin
          port4_object   = port_object_in[5];
          portf_assigned = 1;
        end else if (PRIO_DEPTH[ii*8+:8] > 3 && TX_PORTG_ENABLE && TX_PORTG_PRIORITY == ii && !portg_assigned) begin
          port4_object   = port_object_in[6];
          portg_assigned = 1;
        end else if (PRIO_DEPTH[ii*8+:8] > 3 && TX_PORTH_ENABLE && TX_PORTH_PRIORITY == ii) begin
          port4_object   = port_object_in[7];
        end else begin
          port4_object   = 'hx;
        end


        // fifth port assignment
        if (PRIO_DEPTH[ii*8+:8] > 4 && TX_PORTE_ENABLE && TX_PORTE_PRIORITY == ii && !porte_assigned) begin
          port5_object   = port_object_in[4];
        end else if (PRIO_DEPTH[ii*8+:8] > 4 && TX_PORTF_ENABLE && TX_PORTF_PRIORITY == ii && !portf_assigned) begin
          port5_object   = port_object_in[5];
          portf_assigned = 1;
        end else if (PRIO_DEPTH[ii*8+:8] > 4 && TX_PORTG_ENABLE && TX_PORTG_PRIORITY == ii && !portg_assigned) begin
          port5_object   = port_object_in[6];
          portg_assigned = 1;
        end else if (PRIO_DEPTH[ii*8+:8] > 4 && TX_PORTH_ENABLE && TX_PORTH_PRIORITY == ii) begin
          port5_object   = port_object_in[7];
        end else begin
          port5_object   = 'hx;
        end


        // sixth port assignment
        if (PRIO_DEPTH[ii*8+:8] > 5 && TX_PORTF_ENABLE && TX_PORTF_PRIORITY == ii && !portf_assigned) begin
          port6_object   = port_object_in[5];
        end else if (PRIO_DEPTH[ii*8+:8] > 5 && TX_PORTG_ENABLE && TX_PORTG_PRIORITY == ii && !portg_assigned) begin
          port6_object   = port_object_in[6];
          portg_assigned = 1;
        end else if (PRIO_DEPTH[ii*8+:8] > 5 && TX_PORTH_ENABLE && TX_PORTH_PRIORITY == ii) begin
          port6_object   = port_object_in[7];
        end else begin
          port6_object   = 'hx;
        end


        // seventh port assignment
        if (PRIO_DEPTH[ii*8+:8] > 6 && TX_PORTG_ENABLE && TX_PORTG_PRIORITY == ii && !portg_assigned) begin
          port7_object   = port_object_in[6];
        end else if (PRIO_DEPTH[ii*8+:8] > 6 && TX_PORTH_ENABLE && TX_PORTH_PRIORITY == ii) begin
          port7_object   = port_object_in[7];
        end else begin
          port7_object   = 'hx;
        end


        // eighth port assignment
        if (PRIO_DEPTH[ii*8+:8] > 7 && TX_PORTH_ENABLE && TX_PORTH_PRIORITY == ii) begin
          port8_object   = port_object_in[7];
        end else begin
          port8_object   = 'hx;
        end

      end // end always @*


    // arb_tx_mux priority instance
    srio_gen2_v4_1_16_arb_tx_mux
      #(.TCQ                     (TCQ),
        .TX_ENABLE_FAIRNESS      (TX_ENABLE_FAIRNESS),
        .NUMBER_OF_PORTS         (PRIO_DEPTH[ii*8+:8]))
      arb_tx_mux_inst
       (
        .log_clk                 (log_clk),
        .log_rst_q               (log_rst_q),

        .advance_condition       (advance_condition),

        .LAM_port1_tvalid        (port1_object[0]),
        .LAM_port1_tlast         (port1_object[1]),
        .LAM_port1_tready        (port1_object[2]),
        .LAM_port1_id            (port1_object[TX_OBJECT_WIDTH-1:TX_OBJECT_WIDTH-PORT_ID]),

        .LAM_port2_tvalid        (port2_object[0]),
        .LAM_port2_tlast         (port2_object[1]),
        .LAM_port2_tready        (port2_object[2]),
        .LAM_port2_id            (port2_object[TX_OBJECT_WIDTH-1:TX_OBJECT_WIDTH-PORT_ID]),

        .LAM_port3_tvalid        (port3_object[0]),
        .LAM_port3_tlast         (port3_object[1]),
        .LAM_port3_tready        (port3_object[2]),
        .LAM_port3_id            (port3_object[TX_OBJECT_WIDTH-1:TX_OBJECT_WIDTH-PORT_ID]),

        .LAM_port4_tvalid        (port4_object[0]),
        .LAM_port4_tlast         (port4_object[1]),
        .LAM_port4_tready        (port4_object[2]),
        .LAM_port4_id            (port4_object[TX_OBJECT_WIDTH-1:TX_OBJECT_WIDTH-PORT_ID]),

        .LAM_port5_tvalid        (port5_object[0]),
        .LAM_port5_tlast         (port5_object[1]),
        .LAM_port5_tready        (port5_object[2]),
        .LAM_port5_id            (port5_object[TX_OBJECT_WIDTH-1:TX_OBJECT_WIDTH-PORT_ID]),

        .LAM_port6_tvalid        (port6_object[0]),
        .LAM_port6_tlast         (port6_object[1]),
        .LAM_port6_tready        (port6_object[2]),
        .LAM_port6_id            (port6_object[TX_OBJECT_WIDTH-1:TX_OBJECT_WIDTH-PORT_ID]),

        .LAM_port7_tvalid        (port7_object[0]),
        .LAM_port7_tlast         (port7_object[1]),
        .LAM_port7_tready        (port7_object[2]),
        .LAM_port7_id            (port7_object[TX_OBJECT_WIDTH-1:TX_OBJECT_WIDTH-PORT_ID]),

        .LAM_port8_tvalid        (port8_object[0]),
        .LAM_port8_tlast         (port8_object[1]),
        .LAM_port8_tready        (port8_object[2]),
        .LAM_port8_id            (port8_object[TX_OBJECT_WIDTH-1:TX_OBJECT_WIDTH-PORT_ID]),

        .LAM_port_winner         (port_winner_bus[ii])
       );

    // in case there are no ports of a given priority
    end else                  begin : no_tx_arbiter // if/else generate
      //assign port_winner_bus[ii] = NONE;
      assign port_winner_bus[ii] = PORTA;

    end // if/else generate
  end // for generate
  endgenerate

  // }}} End Priority 0 thru 3 Arbitration -------


  // {{{ Final Arbitration Decision -------
  // higher priority always wins over lower priority
// NOTE CFR - changed to immediate assignment for timing improvement
// Now, there are no other priorities than P1.
  always @* begin
//      if (p3_port_winner != NONE) begin
//        port_winner = p3_port_winner;
//      end else if (p2_port_winner != NONE) begin
//        port_winner = p2_port_winner;
//      end else if (p1_port_winner != NONE) begin
//        port_winner = p1_port_winner;
//      end else if (p0_port_winner != NONE) begin
//        port_winner = p0_port_winner;
//      // default winner
//      end else begin
//        port_winner = NONE;
//      end
      port_winner = p1_port_winner;
  end

  // mux the port winner to the output
  always @* begin
    if (advance_condition) begin
      case (port_winner)
        PORTA   : winning_port_object_d = port_object_in[0];
        PORTB   : winning_port_object_d = port_object_in[1];
        PORTC   : winning_port_object_d = port_object_in[2];
        PORTD   : winning_port_object_d = port_object_in[3];
        PORTE   : winning_port_object_d = port_object_in[4];
        PORTF   : winning_port_object_d = port_object_in[5];
        PORTG   : winning_port_object_d = port_object_in[6];
        //PORTH   : winning_port_object_d = port_object_in[7];
        default : winning_port_object_d = port_object_in[7];
        //default : winning_port_object_d = {'hX,3'h0};
        //default : winning_port_object_d = 0;
        //default : winning_port_object_d = 'hX;
      endcase
    end else begin
      winning_port_object_d = winning_port_object;
    end
  end

  always @(posedge log_clk) begin
//  always @(posedge log_clk or posedge log_rst_q) begin
    if (log_rst_q) begin
      winning_port_object[2:0] <= #TCQ 0;
    end else begin
//    end else if (advance_condition) begin
      winning_port_object[2:0] <= #TCQ winning_port_object_d[2:0];
    end
  end
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      winning_port_object[119:3] <= #TCQ 0;
    end else begin
      winning_port_object[119:3] <= #TCQ winning_port_object_d[119:3];
    end
  end

  // separate the object items into distinct parts
  assign la_lhtx_tdata_pre  = winning_port_object[115:52];
  assign la_lhtx_tkeep_pre  = winning_port_object[51:44];
  assign la_lhtx_tuser_pre  = {winning_port_object[43:10], winning_port_object[3], winning_port_object[8:4]};
  assign la_lhtx_tlast_pre  = winning_port_object[1];
  assign la_lhtx_tvalid_pre = winning_port_object[0] && winning_port_object[2];


  // set the appropriate TREADY signal
  always @* begin
    if (advance_condition) begin
        la_tx_porta_tready_early = 1'b0;
        la_tx_portb_tready_early = 1'b0;
        la_tx_portc_tready_early = 1'b0;
        la_tx_portd_tready_early = 1'b0;
        la_tx_porte_tready_early = 1'b0;
        la_tx_portf_tready_early = 1'b0;
        la_tx_portg_tready_early = 1'b0;
        la_tx_porth_tready_early = 1'b0;
      case (port_winner)
      PORTA   : la_tx_porta_tready_early = port_tvalid_mod[0] && !(la_tx_port_tready_d[0] && ug_tx_port_tlast_q[0]);
      PORTB   : la_tx_portb_tready_early = port_tvalid_mod[1] && !(la_tx_port_tready_d[1] && ug_tx_port_tlast_q[1]);
      PORTC   : la_tx_portc_tready_early = port_tvalid_mod[2] && !(la_tx_port_tready_d[2] && ug_tx_port_tlast_q[2]);
      PORTD   : la_tx_portd_tready_early = port_tvalid_mod[3] && !(la_tx_port_tready_d[3] && ug_tx_port_tlast_q[3]);
      PORTE   : la_tx_porte_tready_early = port_tvalid_mod[4] && !(la_tx_port_tready_d[4] && ug_tx_port_tlast_q[4]);
      PORTF   : la_tx_portf_tready_early = port_tvalid_mod[5] && !(la_tx_port_tready_d[5] && ug_tx_port_tlast_q[5]);
      PORTG   : la_tx_portg_tready_early = port_tvalid_mod[6] && !(la_tx_port_tready_d[6] && ug_tx_port_tlast_q[6]);
      PORTH   : la_tx_porth_tready_early = port_tvalid_mod[7] && !(la_tx_port_tready_d[7] && ug_tx_port_tlast_q[7]);
      default : ;
      endcase
    end else begin
      la_tx_porta_tready_early = la_tx_port_tready_d[0];
      la_tx_portb_tready_early = la_tx_port_tready_d[1];
      la_tx_portc_tready_early = la_tx_port_tready_d[2];
      la_tx_portd_tready_early = la_tx_port_tready_d[3];
      la_tx_porte_tready_early = la_tx_port_tready_d[4];
      la_tx_portf_tready_early = la_tx_port_tready_d[5];
      la_tx_portg_tready_early = la_tx_port_tready_d[6];
      la_tx_porth_tready_early = la_tx_port_tready_d[7];
    end
  end
  always @* begin
    // This is the eval timeout signal, deliberately confusing name
    if (log_packet_first_beat) begin
      la_tx_port_tready_dd[0] = 1'b0;
      la_tx_port_tready_dd[1] = 1'b0;
      la_tx_port_tready_dd[2] = 1'b0;
      la_tx_port_tready_dd[3] = 1'b0;
      la_tx_port_tready_dd[4] = 1'b0;
      la_tx_port_tready_dd[5] = 1'b0;
      la_tx_port_tready_dd[6] = 1'b0;
      la_tx_port_tready_dd[7] = 1'b0;
    end else begin
      la_tx_port_tready_dd[0] = la_tx_porta_tready_early;
      la_tx_port_tready_dd[1] = la_tx_portb_tready_early;
      la_tx_port_tready_dd[2] = la_tx_portc_tready_early;
      la_tx_port_tready_dd[3] = la_tx_portd_tready_early;
      la_tx_port_tready_dd[4] = la_tx_porte_tready_early;
      la_tx_port_tready_dd[5] = la_tx_portf_tready_early;
      la_tx_port_tready_dd[6] = la_tx_portg_tready_early;
      la_tx_port_tready_dd[7] = la_tx_porth_tready_early;
    end
  end
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      la_tx_port_tready_d <= #TCQ 8'h0;
    end else begin
      la_tx_port_tready_d <= #TCQ la_tx_port_tready_dd;
    end
  end

  // }}} End Final Arbitration Decision ---


  // {{{ Pipeline Instantiation -------------------

  assign LA_lhtx_tdata  = la_lhtx_tdata_pre;
  assign LA_lhtx_tkeep  = la_lhtx_tkeep_pre;
  assign LA_lhtx_tuser  = la_lhtx_tuser_pre;
  assign LA_lhtx_tlast  = la_lhtx_tlast_pre;
  assign LA_lhtx_tvalid = la_lhtx_tvalid_pre;
  assign ld_lhtx_tready_pre = LD_lhtx_tready;

//  srio_gen2_v4_1_16_arb_tx_pipe
//    #(.TCQ                    (TCQ))
//    arb_tx_pipe_inst
//    (.log_clk                 (log_clk),
//     .log_rst_q               (log_rst_q),
//
//     .LA_lhtx_tvalid_pre      (la_lhtx_tvalid_pre),
//     .LD_lhtx_tready_pre      (ld_lhtx_tready_pre),
//     .LA_lhtx_tdata_pre       (la_lhtx_tdata_pre),
//     .LA_lhtx_tkeep_pre       (la_lhtx_tkeep_pre),
//     .LA_lhtx_tlast_pre       (la_lhtx_tlast_pre),
//     .LA_lhtx_tuser_pre       (la_lhtx_tuser_pre),
//
//     .LA_lhtx_tvalid          (LA_lhtx_tvalid),
//     .LD_lhtx_tready          (LD_lhtx_tready),
//     .LA_lhtx_tdata           (LA_lhtx_tdata),
//     .LA_lhtx_tkeep           (LA_lhtx_tkeep),
//     .LA_lhtx_tlast           (LA_lhtx_tlast),
//     .LA_lhtx_tuser           (LA_lhtx_tuser)
//   );
  // }}} End of Pipeline Instantiation ------------


  // {{{ Evaluation Core Logic ------------
  // Only generate this is EVAL is set.  This will mask off the incoming valid
  // to be always 0 so no data will be sent out only idles.
  generate if (EVAL) begin : valid_gen
    wire is_valid;

    //The eval logic can not be reset
    srio_gen2_v4_1_16_eval_log_clk  #(
      .TCQ (TCQ)
    ) valid_inst (
      .flag (log_packet_first_beat_d),
      .rst  (1'b0),
      .clk  (log_clk)
     );

  end endgenerate
  always @(posedge log_clk) begin
    if (!EVAL) begin
      log_packet_first_beat <= #TCQ 1'b0;
    end else begin
      log_packet_first_beat <= #TCQ log_packet_first_beat_d;
    end
  end
  // }}} End Evaluation Core Logic --------


  // {{{ Coverage and Assertions ----------

    // *- COVERAGE (cr_LAT_tvalid_coverage)
    // With all ports enabled, cross all combinations of TVALID with ENABLE_FAIRNESS

    // *- COVERAGE (cp_LAT_response_only_request)
    // *- COVERAGE (cp_LAT_response_only_response)
    // Observe the assertion of BT_response_only with and without only a
    // request being queued up.

    // *- COVERAGE (cp_LAT_response_only_mid_packet)
    // Observe BT_response_only assert when in mid_packet, both response and request

    // *- COVERAGE (cp_LAT_response_only_out_of_packet)
    // Observe BT_response_only assert when out of a packet

    // *- COVERAGE (cp_LAT_response_only_on_sof)
    // Observe BT_response_only assert on the same cycle as sof

    // *- COVERAGE (cp_LAT_response_only_on_eof)
    // Observe BT_response_only assert on the same cycle as eof

    // *- COVERAGE (cp_LAT_response_only_alters_tiebreak)
    // Observe BT_response_only assert with a higher priority request and a lower priority
    // response

    // *- COVERAGE (cp_LAT_response_only_single_cycle)
    // Observe BT_response_only assert on a series of single-cycle packets

    // *- COVERAGE (cp_LAT_response_only_cross_tvalid)
    // Observe BT_response_only rise when there is a TVALID on each individual port

    // *- COVERAGE (cp_LAT_maint_only_cross_tvalid)
    // Observe PC_maint_only rise when there is a TVALID on each individual port

    // *- COVERAGE (cp_LAT_stall_sof)
    // Observe a stall on the encoder side on the first beat of a packet

    // *- COVERAGE (cp_LAT_stall_mid)
    // Observe a stall on the encoder side in the middle of the packet

    // *- COVERAGE (cp_LAT_stall_eof)
    // Observe a stall on the encoder side on the last beat of a packet

    // *- COVERAGE (cp_LAT_back_to_back)
    // Observe back-to-back packets with and without ENABLE_FAIRNESS

    // *- COVERAGE (cp_LAT_priority)
    // Observe a higher priority packet when a lower packet is in progress

    // *- COVERAGE (cp_LAT_tvalid_drop_second_beat)
    // Observe TVALID drop on the second beat of a packet

    // *- COVERAGE (cp_LAT_tvalid_drop_mid_packet)
    // Observe TVALID drop mid-packet

    // *- COVERAGE (cp_LAT_tvalid_drop_with_pending_packet)
    // Observe TVALID drop in the middle of a packet, while TVALID of
    // another packet is set

    // *- COVERAGE (cp_LAT_tready_drop_final_beat)
    // Observe TREADY drop on when TLAST asserts

    // *- COVERAGE (cp_LAT_packet_size)
    // Observe incoming packets of sizes 1, 2, 3, and 4+

    // *- COVERAGE (cp_LAT_tvalid_on_tlast)
    // Observe a new, solitary TVALID arrive on TLAST of a packet being serviced

    // *- COVERAGE (cp_LAT_tvalid_1_before_tlast)
    // Observe a new, solitary TVALID arrive one cycle before TLAST of a packet being serviced

    // *- COVERAGE (cp_LAT_tvalid_1_after_tlast)
    // Observe a new, solitary TVALID arrive one cycle after TLAST of a packet being serviced

  // }}} End Coverage and Assertions -------------


endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/log/log_arb/srio_gen2_v4_1_16_eval_log_clk.v#1 $
//----------------------------------------------------------------------
//
// EVAL_LOG_CLK
// Description:
// This is the evaluation timer for the LOG TX which runs on the log_clk
//
// Hierarchy:
// PHY_TOP
//    |___OPLM_TOP
//            |___OPLM_TX
//                    |___EVAL_GT_CLK <-- this module
// ---------------------------------------------------------------------
`timescale 1ps/1ps
// ------------------------------------------------
// below attribute is added to supress the synthesis warnings in vivado tool 8:3332
(* DowngradeIPIdentifiedWarnings="yes" *)
// ------------------------------------------------

module srio_gen2_v4_1_16_eval_log_clk #(
  parameter TCQ     = 100)
(
  output reg  flag  = 0,
  input       rst,
  input       clk
);

  // This clock will operate in the LOG_CLK domain. This module assumes
  // LOG_CLK is running at the highest rate (312.5MHz). It could very well
  // be operating at any frequency. Assuming it runs at the highest rate it
  // guarantees the timeout will not occur before 8 hours, though could trail
  // on for quite a while. However, two other eval timers make certain that
  // full capability won't trail on.
  // 8 hrs -> 480 min -> 28,800 s -> 28,800,000,000 us
  // LOG_CLK (Mhz) | Period (us) | Cycle Count Needed      
  //     312.5     |  .0032      | 9,000,000,000,000 -> (255^5)*8 ~ 7.6

  // Need 5 Stages reguardless of mode (A-E)
  // Initialize all registers to 0 since no reset is attached to this module

  // Stage A
  //------------------------------
  reg   [7:0] a = 0;
  reg         a_out = 0;
  wire        a_ceo;
  wire        a_en;

  assign a_en = 1'b1;

  always @(posedge clk) begin 
    if (rst) begin
      a     <= #TCQ 0;
      a_out <= #TCQ 0;
    end else begin
      if (a_en) begin
        a   <= #TCQ a + 1;
      end
      a_out <= #TCQ a_ceo;
    end
  end

  assign a_ceo = a_en & (&a);

  // Stage B
  //------------------------------
  reg   [7:0] b = 0;
  reg         b_out = 0;
  wire        b_ceo;
  wire        b_en;

  assign b_en = a_out;

  always @(posedge clk) begin
    if (rst) begin
      b     <= #TCQ 0;
      b_out <= #TCQ 0;
    end else begin
      if (b_en) begin
        b   <= #TCQ b + 1;
      end
      b_out <= #TCQ b_ceo;
    end
  end

  assign b_ceo = b_en & (&b);


  // Stage C
  //------------------------------
  reg   [7:0] c = 0;
  reg         c_out = 0;
  wire        c_ceo;
  wire        c_en;

  assign c_en = b_out;

  always @(posedge clk) begin
    if (rst) begin
      c     <= #TCQ 0;
      c_out <= #TCQ 0;
    end else begin
      if (c_en) begin
        c   <= #TCQ c + 1;
      end
      c_out <= #TCQ c_ceo;
    end
  end

  assign c_ceo = c_en & (&c);


  // Stage D
  //------------------------------
  reg   [7:0] d = 0;
  reg         d_out = 0;
  wire        d_ceo;
  wire        d_en;

  assign d_en = c_out;

  always @(posedge clk) begin
    if (rst) begin
      d     <= #TCQ 0;
      d_out <= #TCQ 0;
    end else begin
      if (d_en) begin
        d   <= #TCQ d + 1;
      end
      d_out <= #TCQ d_ceo;
    end
  end

  assign d_ceo = d_en & (&d);


  // Stage E
  //------------------------------
  reg   [7:0] e = 0;
  reg         e_out = 0;
  wire        e_ceo;
  wire        e_en;

  assign e_en = d_out;

  always @(posedge clk) begin
    if (rst) begin
      e     <= #TCQ 0;
      e_out <= #TCQ 0;
    end else begin
      if (e_en) begin
        e   <= #TCQ e + 1;
      end
      e_out <= #TCQ e_ceo;
    end
  end

  assign e_ceo = e_en & (&e);

  // Stage F
  // -----------------------------
  localparam LAST_STAGE_COUNT = 7;
  reg  [3:0]  f = 0;
  wire        f_ceo;
  wire        f_en;

  assign f_en = e_out;

  always @(posedge clk) begin
    if (rst) begin
      f <= #TCQ 0;
    end else begin
      if (f_en) begin
        f <= #TCQ f + 1;
      end
    end
  end

  assign f_ceo = f_en & (f == LAST_STAGE_COUNT);

  // Generate the expire flag
  //------------------------------
  always @(posedge clk) begin
    if (rst) begin
      flag <= #TCQ 0;

    end else if (f_ceo) begin
      flag <= #TCQ 1;
    end
  end

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
//
// ARB_RX
// Description:
// This module holds the transmit logic for the Arbiter
//
// Hierarchy:
// LOG_TOP
//    |_____ARB_TX
//             |_____ARB_TX_USER
//             |_____ARB_TX_MUX
//    |_____ARB_RX
//             |_____ARB_RX_PIPE
// ---------------------------------------------------------------------

`timescale 1ps/1ps

// ------------------------------------------------
// below attribute is added to supress the synthesis warnings in vivado tool 8:3332
(* DowngradeIPIdentifiedWarnings="yes" *)
// ------------------------------------------------

module srio_gen2_v4_1_16_arb_rx_pipe
  #(
   // {{{ Parameter declarations -----------
    parameter TCQ                        = 100,
    parameter DEVICEID_WIDTH             = 8)          // Source/Destination ID width {8,16}
   // }}} ----------------------------------
   (
   // {{{ port declarations ----------------
    // clocks and resets and general signals
    input              log_clk,                  // PHY interface clock
    input              log_rst_q,                // Reset for PHY clock Domain

    // configuration registers
    input       [9:0]  LC_lcsba,                 // Local Configuration Base Address register mask value

    // Header Encoder RX Interface
    input              LE_lhrx_tvalid,           // Valid Packet Beat
    output reg         LA_lhrx_tready,           // Packet Beat Accepted
    input      [63:0]  LE_lhrx_tdata,            // Packet Data
    input       [7:0]  LE_lhrx_tkeep,            // Valid bytes in this beat, only valid on last
    input              LE_lhrx_tlast,            // Last Beat
    input      [39:0]  LE_lhrx_tuser,            // {DEST_ID, SRC_ID, 2'h0, HELLO_FMT, 2'h0, VC, CRF, 1'b0}
    input              LE_unsupported_type,      // The packet has been decoded as an unsupported type

    // Header Encoder RX Interface
    output reg         LE_lhrx_tvalid_q,         // Valid Packet Beat
    input              LA_lhrx_tready_d,         // Packet Beat Accepted
    output reg  [63:0] LE_lhrx_tdata_q,          // Packet Data
    output reg   [7:0] LE_lhrx_tkeep_q,          // Valid bytes in this beat, only valid on last
    output reg         LE_lhrx_tlast_q,          // Last Beat
    output reg  [39:0] LE_lhrx_tuser_q,          // {DEST_ID, SRC_ID, 2'h0, HELLO_FMT, 2'h0, VC, CRF, 1'b0}
    output reg         LE_unsupported_type_q,    // The packet has been decoded as an unsupported type
    output reg  [3:0]  LE_packet_ftype_q,        // Incoming Ftype
    output reg  [3:0]  LE_packet_ttype_q,        // Incoming Ttype
    output reg  [3:0]  LE_packet_stat_q,         // Incoming Stat
    output reg [15:0]  LE_packet_ftype_onehot_q, // one-hot interpretation of ftype
    output reg [15:0]  LE_packet_ttype_onehot_q, // one-hot interpretation of ttype
    output reg [15:0]  LE_packet_stat_onehot_q,  // one-hot interpretation of stat
    output reg  [9:0]  LE_packet_lcsba_q,        // Incoming LCSBA
    output reg         LE_packet_lcsba_hit_q,    // Incoming LCSBA
    output reg         LE_out_of_packet_lhrx_q,  // asserts when the demux is not servicing a packet on lhrx side
    output reg         LE_find_first_beat_q      // used in determining if a packet has begun or not

   // }}} ----------------------------------
   );


  // {{{ local parameters -----------------

  // }}} End local parameters -------------


  // {{{ wire declarations ----------------

  reg   [186:0]   pipeline_in_stg1_d = 0;
  reg   [186:0]   pipeline_in_stg2_d = 0;
  reg   [186:0]   pipeline_in_stg3_d = 0;
  reg   [186:0]   pipeline_in_stg1 = 0;
  reg   [186:0]   pipeline_in_stg2 = 0;
  reg   [186:0]   pipeline_in_stg3 = 0;
  reg             pipeline_vld_stg1, pipeline_vld_stg1_d;
  reg             pipeline_vld_stg2, pipeline_vld_stg2_d;
  reg             pipeline_vld_stg3, pipeline_vld_stg3_d;
  reg     [1:0]   pipeline_in_select, pipeline_in_select_q;

  reg   [3:0]     packet_ftype;                  // Incoming Ftype
  reg   [3:0]     packet_ttype;                  // Incoming Ttype
  reg   [3:0]     packet_stat;                   // Incoming Stat
  reg   [9:0]     packet_lcsba;                  // Incoming LCSBA
  reg             packet_lcsba_hit;              // Hit on LCSBA
  reg   [3:0]     packet_ftype_q;                // Incoming Ftype - registered
  reg   [3:0]     packet_ttype_q;                // Incoming Ttype - registered
  reg   [3:0]     packet_stat_q;                 // Incoming Stat - registered
  reg   [9:0]     packet_lcsba_q;                // Incoming LCSBA - registered
  reg             packet_lcsba_hit_q;            // Hit on LCSBA - registered

  reg             out_of_packet_lhrx;            // asserts when the demux is not servicing a packet on lhrx side
  reg             out_of_packet_lhrx_q;          // asserts when the demux is not servicing a packet on lhrx side
  reg             find_first_beat;               // used in determining if a packet has begun or not

  wire [15:0]     ftype_onehot;
  assign          ftype_onehot[0]  = packet_ftype == 4'h0;
  assign          ftype_onehot[1]  = packet_ftype == 4'h1;
  assign          ftype_onehot[2]  = packet_ftype == 4'h2;
  assign          ftype_onehot[3]  = packet_ftype == 4'h3;
  assign          ftype_onehot[4]  = packet_ftype == 4'h4;
  assign          ftype_onehot[5]  = packet_ftype == 4'h5;
  assign          ftype_onehot[6]  = packet_ftype == 4'h6;
  assign          ftype_onehot[7]  = packet_ftype == 4'h7;
  assign          ftype_onehot[8]  = packet_ftype == 4'h8;
  assign          ftype_onehot[9]  = packet_ftype == 4'h9;
  assign          ftype_onehot[10] = packet_ftype == 4'ha;
  assign          ftype_onehot[11] = packet_ftype == 4'hb;
  assign          ftype_onehot[12] = packet_ftype == 4'hc;
  assign          ftype_onehot[13] = packet_ftype == 4'hd;
  assign          ftype_onehot[14] = packet_ftype == 4'he;
  assign          ftype_onehot[15] = packet_ftype == 4'hf;

  wire [15:0]     ttype_onehot;
  assign          ttype_onehot[0]  = packet_ttype == 4'h0;
  assign          ttype_onehot[1]  = packet_ttype == 4'h1;
  assign          ttype_onehot[2]  = packet_ttype == 4'h2;
  assign          ttype_onehot[3]  = packet_ttype == 4'h3;
  assign          ttype_onehot[4]  = packet_ttype == 4'h4;
  assign          ttype_onehot[5]  = packet_ttype == 4'h5;
  assign          ttype_onehot[6]  = packet_ttype == 4'h6;
  assign          ttype_onehot[7]  = packet_ttype == 4'h7;
  assign          ttype_onehot[8]  = packet_ttype == 4'h8;
  assign          ttype_onehot[9]  = packet_ttype == 4'h9;
  assign          ttype_onehot[10] = packet_ttype == 4'ha;
  assign          ttype_onehot[11] = packet_ttype == 4'hb;
  assign          ttype_onehot[12] = packet_ttype == 4'hc;
  assign          ttype_onehot[13] = packet_ttype == 4'hd;
  assign          ttype_onehot[14] = packet_ttype == 4'he;
  assign          ttype_onehot[15] = packet_ttype == 4'hf;

  wire [15:0]     stat_onehot;
  assign          stat_onehot[0]  = packet_stat == 4'h0;
  assign          stat_onehot[1]  = packet_stat == 4'h1;
  assign          stat_onehot[2]  = packet_stat == 4'h2;
  assign          stat_onehot[3]  = packet_stat == 4'h3;
  assign          stat_onehot[4]  = packet_stat == 4'h4;
  assign          stat_onehot[5]  = packet_stat == 4'h5;
  assign          stat_onehot[6]  = packet_stat == 4'h6;
  assign          stat_onehot[7]  = packet_stat == 4'h7;
  assign          stat_onehot[8]  = packet_stat == 4'h8;
  assign          stat_onehot[9]  = packet_stat == 4'h9;
  assign          stat_onehot[10] = packet_stat == 4'ha;
  assign          stat_onehot[11] = packet_stat == 4'hb;
  assign          stat_onehot[12] = packet_stat == 4'hc;
  assign          stat_onehot[13] = packet_stat == 4'hd;
  assign          stat_onehot[14] = packet_stat == 4'he;
  assign          stat_onehot[15] = packet_stat == 4'hf;


  // }}} End wire declarations ------------


  // {{{ Receive Path Pipeline ------------
  always @* begin
    pipeline_in_stg1_d = pipeline_in_stg1;
    if (LE_lhrx_tvalid && LA_lhrx_tready) begin
      pipeline_in_stg1_d = {packet_lcsba_hit, ftype_onehot, ttype_onehot, stat_onehot, out_of_packet_lhrx,
                           find_first_beat, packet_ftype, packet_ttype, packet_stat, packet_lcsba,
                           LE_unsupported_type, LE_lhrx_tlast, LE_lhrx_tkeep, LE_lhrx_tuser, LE_lhrx_tdata};
    end

    pipeline_in_stg2_d = pipeline_in_stg2;
    if ((!pipeline_vld_stg2 || !pipeline_vld_stg3) || (LE_lhrx_tvalid_q && LA_lhrx_tready_d)) begin
      pipeline_in_stg2_d = pipeline_in_stg1;
    end

    pipeline_in_stg3_d = pipeline_in_stg3;
    if ((!pipeline_vld_stg3) || (LE_lhrx_tvalid_q && LA_lhrx_tready_d)) begin
      pipeline_in_stg3_d = pipeline_in_stg2;
    end
  end

  always @(posedge log_clk) begin
    if (log_rst_q) begin
      pipeline_in_stg1 <= #TCQ 1'b0;
      pipeline_in_stg2 <= #TCQ 1'b0;
      pipeline_in_stg3 <= #TCQ 1'b0;
    end else begin
      pipeline_in_stg1 <= #TCQ pipeline_in_stg1_d;
      pipeline_in_stg2 <= #TCQ pipeline_in_stg2_d;
      pipeline_in_stg3 <= #TCQ pipeline_in_stg3_d;
    end
  end

  always @* begin
    pipeline_vld_stg1_d = pipeline_vld_stg1;
    if (LE_lhrx_tvalid && LA_lhrx_tready) begin
      pipeline_vld_stg1_d = 1'b1;
    end else if (!pipeline_vld_stg2 || !pipeline_vld_stg3) begin
      pipeline_vld_stg1_d = 1'b0;
    end else if (LE_lhrx_tvalid_q && LA_lhrx_tready_d) begin
      pipeline_vld_stg1_d = 1'b0;
    end

    pipeline_vld_stg2_d = pipeline_vld_stg2;
    if (pipeline_vld_stg1) begin
      pipeline_vld_stg2_d = !((pipeline_in_select_q == 2'b01) && (LE_lhrx_tvalid_q && LA_lhrx_tready_d));
    end else if (!pipeline_vld_stg3 || (pipeline_in_select_q == 2'b11 || pipeline_in_select_q == 2'b10) &&
                  (LE_lhrx_tvalid_q && LA_lhrx_tready_d)) begin
      pipeline_vld_stg2_d = 1'b0;
    end

    pipeline_vld_stg3_d = pipeline_vld_stg3;
    if (pipeline_vld_stg2) begin
      pipeline_vld_stg3_d = !((pipeline_in_select_q == 2'b10) && (LE_lhrx_tvalid_q && LA_lhrx_tready_d));
    end else if (pipeline_in_select_q == 2'b11 && (LE_lhrx_tvalid_q && LA_lhrx_tready_d)) begin
      pipeline_vld_stg3_d = 1'b0;
    end
  end

  always @(posedge log_clk) begin
    if (log_rst_q) begin
      pipeline_vld_stg1 <= #TCQ 1'b0;
      pipeline_vld_stg2 <= #TCQ 1'b0;
      pipeline_vld_stg3 <= #TCQ 1'b0;
    end else begin
      pipeline_vld_stg1 <= #TCQ pipeline_vld_stg1_d;
      pipeline_vld_stg2 <= #TCQ pipeline_vld_stg2_d;
      pipeline_vld_stg3 <= #TCQ pipeline_vld_stg3_d;
    end
  end

  always @* begin
    casex ({pipeline_vld_stg3_d, pipeline_vld_stg2_d, pipeline_vld_stg1_d})
      3'b1xx  : pipeline_in_select = 2'b11;
      3'b01x  : pipeline_in_select = 2'b10;
      3'b001  : pipeline_in_select = 2'b01;
      default : pipeline_in_select = 2'b00;
    endcase
  end
  always @(posedge log_clk) begin
    pipeline_in_select_q <= #TCQ pipeline_in_select;
  end
  // }}} End Receive Path Pipeline --------


  // {{{ Packet Decode Logic --------------

  // determine when out-of-packet in order to find the first beat of the next packet
  // This is done pre-pipeline in order to reduce the number of logic levels on the demux

  always @* begin
    out_of_packet_lhrx = out_of_packet_lhrx_q;
    if (LA_lhrx_tready && LE_lhrx_tvalid && LE_lhrx_tlast) begin
      out_of_packet_lhrx = 1'b1;
    end else if (LE_lhrx_tvalid) begin
      out_of_packet_lhrx = 1'b0;
    end
  end
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      out_of_packet_lhrx_q           <= #TCQ 1'b1;
    end else begin
      out_of_packet_lhrx_q           <= #TCQ out_of_packet_lhrx;
    end
  end

  // For decoding the packet details - FTYPE, TTYPE, STAT:
  // asserts when looking for the first beat of data on the LHRX side
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      find_first_beat <= #TCQ 1'b1;
    end else if (out_of_packet_lhrx) begin
      find_first_beat <= #TCQ 1'b1;
    end else if (LA_lhrx_tready && LE_lhrx_tvalid) begin
      find_first_beat <= #TCQ 1'b0;
    end
  end

  // decode the appropriate fields - FTYPE, TTYPE, STAT
  always @* begin
    packet_ftype     = packet_ftype_q;
    packet_ttype     = packet_ttype_q;
    packet_stat      = packet_stat_q;
    packet_lcsba     = packet_lcsba_q;
    packet_lcsba_hit = packet_lcsba_hit_q;
    if (find_first_beat) begin
      // HELLO Format in use:
      if (LE_lhrx_tuser[5]) begin
        packet_ftype     = LE_lhrx_tdata[55:52];
        packet_ttype     = LE_lhrx_tdata[51:48];
        packet_stat      = LE_lhrx_tdata[35] == 0 ? 4'h0 : 4'h7;
        packet_lcsba     = LE_lhrx_tdata[33:24];
        packet_lcsba_hit = LE_lhrx_tdata[33:24] == LC_lcsba;
      // Native sRIO in use:
      end else begin
        packet_ftype     = LE_lhrx_tdata[3:0];
        packet_ttype     = DEVICEID_WIDTH == 16 ? LE_lhrx_tdata[47:44] : LE_lhrx_tdata[31:28];
        packet_stat      = DEVICEID_WIDTH == 16 ? LE_lhrx_tdata[43:40] : LE_lhrx_tdata[27:24];
        packet_lcsba     = 10'h0; // not supported for Native sRIO
        packet_lcsba_hit = 1'b0;
      end
    end
  end
  always @(posedge log_clk) begin
    packet_ftype_q     <= #TCQ packet_ftype;
    packet_ttype_q     <= #TCQ packet_ttype;
    packet_stat_q      <= #TCQ packet_stat;
    packet_lcsba_q     <= #TCQ packet_lcsba;
    packet_lcsba_hit_q <= #TCQ packet_lcsba_hit;
  end

  // }}} End of Packet Decode Logic -------


  // {{{ Assignments to Ports -------------
  wire         LE_unsupported_type_int    = pipeline_in_select == 2'b11 ? pipeline_in_stg3_d[113] :
                                      pipeline_in_select == 2'b10 ? pipeline_in_stg2_d[113] :
                                                                    pipeline_in_stg1_d[113];
  wire         LE_lhrx_tlast_int          = pipeline_in_select == 2'b11 ? pipeline_in_stg3_d[112] :
                                      pipeline_in_select == 2'b10 ? pipeline_in_stg2_d[112] :
                                                                    pipeline_in_stg1_d[112];
  wire [63:0]  LE_lhrx_tdata_int          = pipeline_in_select == 2'b11 ? pipeline_in_stg3_d[63:0] :
                                      pipeline_in_select == 2'b10 ? pipeline_in_stg2_d[63:0] :
                                                                    pipeline_in_stg1_d[63:0];
  wire  [7:0]  LE_lhrx_tkeep_int          = pipeline_in_select == 2'b11 ? pipeline_in_stg3_d[111:104] :
                                      pipeline_in_select == 2'b10 ? pipeline_in_stg2_d[111:104] :
                                                                    pipeline_in_stg1_d[111:104];
  wire [39:0]  LE_lhrx_tuser_int          = pipeline_in_select == 2'b11 ? pipeline_in_stg3_d[103:64] :
                                      pipeline_in_select == 2'b10 ? pipeline_in_stg2_d[103:64] :
                                                                    pipeline_in_stg1_d[103:64];

  wire  [3:0]  LE_packet_ftype_int        = pipeline_in_select == 2'b11 ? pipeline_in_stg3_d[135:132] :
                                      pipeline_in_select == 2'b10 ? pipeline_in_stg2_d[135:132] :
                                                                    pipeline_in_stg1_d[135:132];
  wire  [3:0]  LE_packet_ttype_int        = pipeline_in_select == 2'b11 ? pipeline_in_stg3_d[131:128] :
                                      pipeline_in_select == 2'b10 ? pipeline_in_stg2_d[131:128] :
                                                                    pipeline_in_stg1_d[131:128];
  wire  [3:0]  LE_packet_stat_int         = pipeline_in_select == 2'b11 ? pipeline_in_stg3_d[127:124] :
                                      pipeline_in_select == 2'b10 ? pipeline_in_stg2_d[127:124] :
                                                                    pipeline_in_stg1_d[127:124];
  wire  [9:0]  LE_packet_lcsba_int        = pipeline_in_select == 2'b11 ? pipeline_in_stg3_d[123:114] :
                                      pipeline_in_select == 2'b10 ? pipeline_in_stg2_d[123:114] :
                                                                    pipeline_in_stg1_d[123:114];
  wire         LE_out_of_packet_lhrx_int  = pipeline_in_select == 2'b11 ? pipeline_in_stg3_d[137] :
                                      pipeline_in_select == 2'b10 ? pipeline_in_stg2_d[137] :
                                                                    pipeline_in_stg1_d[137];
  wire         LE_find_first_beat_int     = pipeline_in_select == 2'b11 ? pipeline_in_stg3_d[136] :
                                      pipeline_in_select == 2'b10 ? pipeline_in_stg2_d[136] :
                                                                    pipeline_in_stg1_d[136];

  wire [15:0]  LE_packet_stat_onehot_int  = pipeline_in_select == 2'b11 ? pipeline_in_stg3_d[153:138] :
                                      pipeline_in_select == 2'b10 ? pipeline_in_stg2_d[153:138] :
                                                                    pipeline_in_stg1_d[153:138];
  wire [15:0]  LE_packet_ttype_onehot_int = pipeline_in_select == 2'b11 ? pipeline_in_stg3_d[169:154] :
                                      pipeline_in_select == 2'b10 ? pipeline_in_stg2_d[169:154] :
                                                                    pipeline_in_stg1_d[169:154];
  wire [15:0]  LE_packet_ftype_onehot_int = pipeline_in_select == 2'b11 ? pipeline_in_stg3_d[185:170] :
                                      pipeline_in_select == 2'b10 ? pipeline_in_stg2_d[185:170] :
                                                                    pipeline_in_stg1_d[185:170];
  wire         LE_packet_lcsba_hit_int    = pipeline_in_select == 2'b11 ? pipeline_in_stg3_d[186] :
                                      pipeline_in_select == 2'b10 ? pipeline_in_stg2_d[186] :
                                                                    pipeline_in_stg1_d[186];


  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LE_lhrx_tvalid_q <= #TCQ 1'b0;
      LA_lhrx_tready   <= #TCQ 1'b0;
    end else begin
      LE_lhrx_tvalid_q <= #TCQ pipeline_vld_stg3_d || pipeline_vld_stg2_d || pipeline_vld_stg1_d;
      LA_lhrx_tready   <= #TCQ !(pipeline_vld_stg3_d && pipeline_vld_stg2_d && pipeline_vld_stg1_d);
    end
  end

  always @(posedge log_clk) begin
    LE_unsupported_type_q    <= #TCQ LE_unsupported_type_int;
    LE_lhrx_tlast_q          <= #TCQ LE_lhrx_tlast_int;
    LE_lhrx_tdata_q          <= #TCQ LE_lhrx_tdata_int;
    LE_lhrx_tkeep_q          <= #TCQ LE_lhrx_tkeep_int;
    LE_lhrx_tuser_q          <= #TCQ LE_lhrx_tuser_int;
    LE_packet_ftype_q        <= #TCQ LE_packet_ftype_int;
    LE_packet_ttype_q        <= #TCQ LE_packet_ttype_int;
    LE_packet_stat_q         <= #TCQ LE_packet_stat_int;
    LE_packet_lcsba_q        <= #TCQ LE_packet_lcsba_int;
    LE_out_of_packet_lhrx_q  <= #TCQ LE_out_of_packet_lhrx_int;
    LE_find_first_beat_q     <= #TCQ LE_find_first_beat_int;
    LE_packet_stat_onehot_q  <= #TCQ LE_packet_stat_onehot_int;
    LE_packet_ttype_onehot_q <= #TCQ LE_packet_ttype_onehot_int;
    LE_packet_ftype_onehot_q <= #TCQ LE_packet_ftype_onehot_int;
    LE_packet_lcsba_hit_q    <= #TCQ LE_packet_lcsba_hit_int;
  end

  // }}} End Assignments to Ports ---------


endmodule
// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/log/log_hello/srio_gen2_v4_1_16_hello_encoder.v#1 $
//----------------------------------------------------------------------
//
// HELLO_ENCODER
// Description:
// This module converts packets from Buffer Native format to sRIO Native
// or HELLO format based on FTYPE. It sits in the LOG RX data path
// between the RX Buffer and the LOG RX Arbiter.
//
// Hierarchy:
// LOG_TOP
//    |___HELLO_ENCODER - this module
// ---------------------------------------------------------------------

`timescale 1ps/1ps

module srio_gen2_v4_1_16_hello_encoder
#(
  parameter TCQ               = 100, // in ps
  parameter DEVICEID_WIDTH    =   8, // Indicates Source/Dest ID width {8, 16}
  parameter TARGET_NREAD      =   1, // If 1, core may sink NRead transactions {0, 1}
  parameter TARGET_NWRITE     =   1, // If 1, core may sink NWrite transactions {0, 1}
  parameter TARGET_NWRITE_R   =   1, // If 1, core may sink NWrite_R transactions {0, 1}
  parameter TARGET_SWRITE     =   1, // If 1, core may sink SWrite transactions {0, 1}
  parameter TARGET_DB         =   1, // If 1, core may sink Doorbell transactions {0, 1}
  parameter TARGET_DS         =   1, // If 1, core may sink Data Streaming {0, 1}
  parameter TARGET_ATOMIC     =   1, // If 1, core may sink Atomic transactions {0, 1}
  parameter INIT_NREAD        =   1, // If 1, core may initiate NRead transactions {0, 1}
  parameter INIT_NWRITE_R     =   1, // If 1, core may initiate NWrite_R transactions {0, 1}
  parameter INIT_DB           =   1, // If 1, core may initiate Doorbell transactions {0, 1}
  parameter INIT_ATOMIC       =   1, // If 1, core may initiate Atomic transactions {0, 1}
  parameter MSG_SINK_SINGLE   =   1, // If 1, core may sink single segment msg transactions {0, 1}
  parameter MSG_SINK_MULTI    =   1, // If 1, core may sink multi-segment msg transactions {0, 1}
  parameter MSG_INIT_SINGLE   =   1, // If 1, core may initiate single segment msg transactions {0, 1}
  parameter MSG_INIT_MULTI    =   1, // If 1, core may initiate multi-segment msg transactions {0, 1}
  parameter PORT_IO_HELLO     =   1, // The I/O Port uses HELLO format {0,1}
  parameter PORT_MSG_HELLO    =   1, // The Messaging Port uses HELLO format {0,1}
  parameter PORT_MAINT_HELLO  =   1) // The Maintenance Port uses HELLO format {0,1}
(
  // {{{ Port Declarations
  // System Signals
  input                         log_clk,
  input                         log_rst,

  // RX Buffer Interface
  input                         BR_bufr_tvalid,         // Valid packet beat
  output                        LE_bufr_tready,         // Packet beat accepted
  input      [63:0]             BR_bufr_tdata,          // Packet data
  input      [7:0]              BR_bufr_tkeep,          // Valid bytes in this beat, only valid on last
  input                         BR_bufr_tlast,          // Last beat
  input      [7:0]              BR_bufr_tuser,          // {5'h00, VC, CRF, 1'b0}

  // LOG Arbiter Interface
  output reg                    LE_lhrx_tvalid,         // Valid packet beat
  input                         LA_lhrx_tready,         // Packet beat accepted
  output reg [63:0]             LE_lhrx_tdata = 0,      // Packet data
  output reg [7:0]              LE_lhrx_tkeep = 8'hFF,  // Valid bytes in this beat, only valid on last
  output reg                    LE_lhrx_tlast = 0,      // Last beat
  output reg [39:0]             LE_lhrx_tuser = 0,      // {SrcID, DestID, 5'h00, VC, CRF, 1'b0}
  output reg                    LE_unsupported_type     // The packet has been decoded as an unsupported type
  // }}} end Port Declarations
);

  // {{{ Local Parameters

  // Spec defined parameters
  // ------------------------------------------------------------

  //  + {{{ Transactions to encode +
  localparam ENCODE_NREAD           = PORT_IO_HELLO    && TARGET_NREAD;
  localparam ENCODE_NREADATOMIC     = PORT_IO_HELLO    && TARGET_ATOMIC;
  localparam ENCODE_NWRITE          = PORT_IO_HELLO    && TARGET_NWRITE;
  localparam ENCODE_NWRITE_R        = PORT_IO_HELLO    && TARGET_NWRITE_R;
  localparam ENCODE_NWRITEATOMIC    = PORT_IO_HELLO    && TARGET_ATOMIC;
  localparam ENCODE_SWRITE          = PORT_IO_HELLO    && TARGET_SWRITE;
  localparam ENCODE_MAINT           = PORT_MAINT_HELLO;
  localparam ENCODE_DB              = PORT_IO_HELLO    && TARGET_DB;
  localparam ENCODE_DS              = PORT_IO_HELLO    && TARGET_DS;
  localparam ENCODE_MSG             = PORT_MSG_HELLO   && (MSG_SINK_SINGLE || MSG_SINK_MULTI);
  localparam ENCODE_RESPWDATA       = PORT_IO_HELLO    && (INIT_NREAD || INIT_ATOMIC);
  localparam ENCODE_RESPNODATA      = PORT_IO_HELLO    && (INIT_DB || INIT_NWRITE_R);
  localparam ENCODE_RESPMSG         = PORT_MSG_HELLO   && (MSG_INIT_SINGLE || MSG_INIT_MULTI);
  //  + }}} Transactions to encode  +

  // Ftypes of RapidIO spec-defined packet types
  localparam [3:0] FTYPE_NREAD      = 4'b0010;
  localparam [3:0] FTYPE_NWRITE     = 4'b0101;
  localparam [3:0] FTYPE_SWRITE     = 4'b0110;
  localparam [3:0] FTYPE_MAINT      = 4'b1000;
  localparam [3:0] FTYPE_DS         = 4'b1001;
  localparam [3:0] FTYPE_DB         = 4'b1010;
  localparam [3:0] FTYPE_MSG        = 4'b1011;
  localparam [3:0] FTYPE_RESP       = 4'b1101;

  // Parameters used just in this module
  // ------------------------------------------------------------
  localparam HADDR_WIDTH = (DEVICEID_WIDTH == 8) ? 24 : 8; // Width of high address (number of address bits on first DWORD)
  localparam LADDR_WIDTH = 29 - HADDR_WIDTH;               // Width of low address (number of address bits on second DWORD)
  // Short (<1 DWORD) headers are for FTYPEs 11 and 13 (plus 6 and 10 if using 8-bit device IDs)
  localparam SHORT_HEADERS_ONLY = ((!ENCODE_SWRITE && !ENCODE_DB && !ENCODE_DS) || (DEVICEID_WIDTH == 8 )) &&
                                    !ENCODE_NREAD  && !ENCODE_NREADATOMIC && !ENCODE_MAINT   &&
                                    !ENCODE_NWRITE && !ENCODE_NWRITE_R    && !ENCODE_NWRITEATOMIC;
  // Long (>1 DWORD) headers are for FTYPEs 2, 5, and 8 (plus 6 and 10 if using 16-bit device IDs)
  localparam LONG_HEADERS_ONLY =  ((!ENCODE_SWRITE && !ENCODE_DB && !ENCODE_DS) || (DEVICEID_WIDTH == 16)) &&
                                    !ENCODE_MSG    && !ENCODE_RESPWDATA   && !ENCODE_RESPNODATA && !ENCODE_RESPMSG;
  // }}} end Local Parameters


  // {{{ Wire Declarations
  reg                     log_rst_q = 1;

  reg  [7:0]              bufr_keep = 0;  // Registered verison of BR_bufr_tkeep
  reg  [63:0]             bufr_data = 0;  // Registered verison of BR_bufr_tdata
  reg  [7:0]              bufr_user = 0;  // Registered verison of BR_bufr_tuser
  reg                     bufr_last = 0;  // Registered verison of BR_bufr_tlast
  reg                     bufr_last_q = 0;  // Registered verison of BR_bufr_tlast
  reg                     bufr_sof  = 0;  // The data on bufr_data is the sof
  reg                     bufr_valid;     // Registered verison of BR_bufr_tvalid
  wire                    bufr_active_d;  // New valid data on BR_bufr_data (LE_bufr_ready && BR_bufr_valid)
  reg                     bufr_active;    // registered version of bufr_active_d
  wire [63:0]             srio_data;      // Un-swizzled verison of bufr_data
  wire [7:0]              srio_tkeep;      // Un-swizzled verison of bufr_tkeep
  // FIXME CFR - don't want to remove until I know I'm right
  //reg                     bufr_last_hold; // BR_bufr_tlast captured on bufr_active_d, used to create sof
  reg                     bufr_sof_hold;  // bufr_last_hold captured on bufr_active_d, used to identify second beat
  // FIXME CFR - don't want to remove until I know I'm right
  //wire                    bufr_first;     // The data on bufr_data is the first beat of the packet
  wire                    bufr_second;    // The data on bufr_data is the second beat of the packet
  wire                    arb_stall;      // The arbiter is stalling (deasserting ready while valid data present)
  reg                     arb_stall_q;    // Registered version of arb_stall
  reg                     arb_stall_vld;  // Indicate whether there's valid data in the pipe coming out of a stall
  reg                     arb_stall_sof;  // Indicate whether there was an sof at the time of the stall

  // Fields valid on bufr_sof use *_bt1 naming convention
  wire                    crf_bt1;        // CRF of rcvd packet, valid on bufr_sof
  wire [1:0]              prio_bt1;       // Priority of rcvd packet, valid on bufr_sof
  wire [3:0]              ftype_bt1;      // FTYPE of rcvd packet, valid on bufr_sof
  wire [15:0]             destid_bt1;     // Destination ID of rcvd packet, valid on bufr_sof
  wire [15:0]             srcid_bt1;      // Source ID of rcvd packet, valid on bufr_sof
  wire [3:0]              ttype_bt1;      // TTYPE of rcvd packet, valid on bufr_sof
  wire [3:0]              sizestat_bt1;   // Size/Status of rcvd packet, valid on bufr_sof
  reg  [3:0]              sizestat_bt2;   // Size/Status of rcvd packet, valid on bufr_sof
  wire [7:0]              tid_bt1;        // TID of rcvd packet, valid on bufr_sof
  wire [HADDR_WIDTH-1:0]  haddr_bt1;      // The high portion of address on the rcvd packet, valid on bufr_sof
  wire                    ok_bt1;         // Interpretation of status of rcvd packet, valid on bufr_sof
  wire [33:0]             swr_addr_bt1;   // The address of a rcvd SWRITE, valid on bufr_sof
  wire [3:0]              msglen_bt1;     // MSGLEN of rcvd packet, valid on bufr_sof for msg packet
  wire [1:0]              letter_bt1;     // LETTER of rcvd packet, valid on bufr_sof for msg packet
  wire [1:0]              mbox_bt1;       // MBOX of rcvd packet, valid on bufr_sof for msg packet
  wire [3:0]              msgseg_bt1;     // MSGSEG of rcvd packet, valid on bufr_sof for msg packet
  wire [3:0]              xmbox_bt1;      // XMBOX of rcvd packet, valid on bufr_sof for msg packet
  reg                     bad_ssize;      // A bad ssize was decoded from sizestat
  reg  [7:0]              ssize_bt1;      // SSIZE of rcvd packet, valid on bufr_sof for msg packet

  // Fields valid on bufr_second use *_bt2 naming convention
  reg                     crf_bt2;        // CRF of rcvd packet, valid on bufr_second
  reg  [1:0]              prio_bt2;       // Priority of rcvd packet, valid on bufr_second
  reg  [3:0]              ttype_bt2;      // TTYPE of rcvd packet, valid on bufr_second
  reg  [3:0]              rdwrsize_bt2;   // RDSIZE/WRSIZE of rcvd packet, valid on bufr_second
  reg  [7:0]              tid_bt2;        // TID of rcvd packet, valid on bufr_second
  reg  [HADDR_WIDTH-1:0]  haddr_bt2;      // High address bits of rcvd packet, valid on bufr_second
  reg                     ok_bt2;         // Interpretation of status of rcvd packet, valid on bufr_second
  reg  [23:0]             swr_haddr_bt2;  // The high address bits for an SWRITE, valid on bufr_second
  wire [33:0]             swr_addr_bt2;   // Address for 16-bit device ID mode SWRITE, valid on bufr_second
  wire [LADDR_WIDTH-1:0]  laddr_bt2;      // Low address bits of rcvd packet, valid on bufr_second
  wire                    wdptr_bt2;      // WDPTR of rcvd packet, valid on bufr_second
  wire [1:0]              xamsbs_bt2;     // XAMSBS of rcvd packet, valid on bufr_second
  reg                     bad_rdwrsize;   // The decode of rdsize/wrsize and wdptr did not find a valid combo
  reg  [2:0]              addr_lsb_bt2;   // The lower address bits for the HELLO formatted packet
  reg  [7:0]              hello_size_bt2; // The size for the HELLO formatted packet
  wire [7:0]              maint_size_bt2; // The size for a maintenance packet (masked to 0's for MRESPs)
  wire [33:0]             addr_bt2;       // The full HELLO address, valid on bufr_second
  reg  [3:0]              ftype_hold = 0; // The FTYPE captured on SOF so that it's available throughout the pkt
  reg  [3:0]              ttype_hold = 0; // The TTYPE captured on SOF so that it's available throughout the pkt
  wire [3:0]              bufr_ftype;     // The FTYPE of the packet on the bufr interface, valid throughout the pkt
  wire [3:0]              bufr_ttype;     // The TTYPE of the packet on the bufr interface, valid throughout the pkt
  reg  [55:0]             srio_data_hold; // srio_data registered on bufr_active_d, used for data alignment
  reg  [7:0]              srio_tkeep_hold; // srio_tkeep registered on bufr_active_d, used for data alignment
  reg                     hello_encode;   // The pkt will be encoded as HELLO (else will be passed in sRIO Native)
  reg                     hello_encode_q; // Registered version of hello_encode used after sof to ease timing
  reg                     unsupported_type_d; // The packet has an unsupported FTYPE/TTYPE (including user-def)
  reg                     header_stage;   // The HELLO encoder is forming the header beat
  reg                     data_stage;     // The HELLO encoder is forming a data beat
  reg  [63:0]             hello_header;   // The HELLO formatted header field, valid on header_stage
  reg  [63:0]             hello_data;     // The aligned data for the HELLO packet, valid on data_stage
  reg  [7:0]              hello_tkeep;     // The aligned data for the HELLO packet, valid on data_stage
  wire                    long_header_ftype9; 
  wire                    short_header_ftype9; 
  wire                    pkt_extend_d;
  // }}} end Wire Declarations




  // {{{ Register Reset
  // Register the reset before use to minimize fanout
  always @(posedge log_clk) begin
    log_rst_q         <= #TCQ log_rst;
  end
  // }}} end Register Reset

  // {{{ Register Core Inputs

  // IPCV - Using BR_bufr_tvalid unregistered
  assign bufr_active_d = BR_bufr_tvalid && LE_bufr_tready; // bufr interface is active when ready && valid

  // Register the bufr_active_d signal to know when the data registered from the interface is fresh
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      bufr_active    <= #TCQ 1'b0;
      bufr_last_q    <= #TCQ 1'b0;
    end else begin
      bufr_active    <= #TCQ bufr_active_d;
      bufr_last_q    <= #TCQ bufr_last;
    end
  end

  // Register core inputs as recommended in IP Checklist
  always @(posedge log_clk) begin
    // No reset to reduce fanout - Not needed because data signals are only sampled on valid cycles
    if (bufr_active_d || pkt_extend_d) begin
      bufr_keep     <= #TCQ BR_bufr_tkeep;
      bufr_data     <= #TCQ BR_bufr_tdata;
      bufr_user     <= #TCQ BR_bufr_tuser;
      bufr_last     <= #TCQ BR_bufr_tlast;
      if (bufr_active_d)
      bufr_sof      <= #TCQ BR_bufr_tuser[3]&& BR_bufr_tkeep[3];
    end else if (!arb_stall) begin
      bufr_last     <= #TCQ 1'b0;
      bufr_sof      <= #TCQ 1'b0;
    end
  end

  // Un-swizzle the data (convert from Buffer Native format to sRIO Native) for easier header parsing
  assign srio_data    = {bufr_data[7:0],  bufr_data[15:8], bufr_data[23:16],bufr_data[31:24],
                         bufr_data[39:32],bufr_data[47:40],bufr_data[55:48],bufr_data[63:56]};

  assign srio_tkeep =  {bufr_keep[0],bufr_keep[1],bufr_keep[2],bufr_keep[3],bufr_keep[4],bufr_keep[5],bufr_keep[6],bufr_keep[7]};

  // Register the data so that it can be shifted onto the next byte as needed
  always @(posedge log_clk) begin
    // No reset needed because only sampled when data is valid
    if (((bufr_active_d || bufr_active)&& !arb_stall) || (arb_stall_q && !arb_stall && arb_stall_vld)) begin
      srio_data_hold   <= #TCQ srio_data[55:0];
      srio_tkeep_hold   <= #TCQ srio_tkeep;
    end
  end

  // }}} end Register Core Inputs

  // {{{ Create Control Signals

  // Keep track of first and second beat of data
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      // FIXME CFR - don't want to remove until I know I'm right
      //bufr_last_hold  <= #TCQ 1'b1; // Reset to one so that sof asserts for the first frame
      bufr_sof_hold   <= #TCQ 1'b0;
    end else if (bufr_active) begin
      // FIXME CFR - don't want to remove until I know I'm right
      //bufr_last_hold  <= #TCQ bufr_last;
      bufr_sof_hold   <= #TCQ bufr_sof && !bufr_last;
    end
  end

  // Set flags to keep track of the first and second beats of data on the bufr registers
  // FIXME CFR - don't want to remove until I know I'm right
  //assign bufr_first  = bufr_active && bufr_last_hold;
  assign bufr_second = bufr_active && bufr_sof_hold;

  // Check for a stall by the arbiter (when there is valid data but the arb does not accept it)
  assign arb_stall = LE_lhrx_tvalid && !LA_lhrx_tready;

  // Register the arbiter stall flag to use to find the falling edge
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      arb_stall_q     <= #TCQ 1'b0;
    end else begin
      arb_stall_q     <= #TCQ arb_stall;
    end
  end

  // Keep track of whether there's valid data in the pipe when the arb stall releases
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      arb_stall_vld   <= #TCQ 1'b0;
      arb_stall_sof   <= #TCQ 1'b0;
    end else if (arb_stall && !arb_stall_q) begin
      arb_stall_vld   <= #TCQ (!hello_encode && bufr_active) || header_stage || data_stage;
      arb_stall_sof   <= #TCQ bufr_sof;
    end
  end

  // Determine sof on bufr/srio_data buses
  // FIXME CFR - don't want to remove until I know I'm right
  //assign bufr_sof = bufr_first || ((!arb_stall && arb_stall_q) && arb_stall_sof);

  // }}} end Create Control Signals

  // {{{ Parse Received Packet

  // Decode first-beat header fields
  // I/O Fields
  assign crf_bt1      = bufr_user[1];
  assign prio_bt1     = srio_data[63:62];
  assign ftype_bt1    = srio_data[59:56];
  assign destid_bt1   = (DEVICEID_WIDTH == 8) ? {8'b0,srio_data[55:48]} : srio_data[55:40];
  assign srcid_bt1    = (DEVICEID_WIDTH == 8) ? {8'b0,srio_data[47:40]} : srio_data[39:24];
  assign ttype_bt1    = (DEVICEID_WIDTH == 8) ? srio_data[39:36] : srio_data[23:20];
  assign sizestat_bt1 = (DEVICEID_WIDTH == 8) ? srio_data[35:32] : srio_data[19:16];
  assign tid_bt1      = (DEVICEID_WIDTH == 8) ? srio_data[31:24] : srio_data[15:8];
  assign haddr_bt1    = (DEVICEID_WIDTH == 8) ? srio_data[23:0]  : srio_data[7:0];
  assign ok_bt1       = (({1'b0,ftype_bt1} == FTYPE_RESP[3:0]) ||
                        (({1'b0,ftype_bt1} == FTYPE_MAINT[3:0]) && ttype_bt1[1])) ?
                         (sizestat_bt1 == 4'h0) : 1'b1;   // Set to one unless response
  assign swr_addr_bt1 = (DEVICEID_WIDTH == 8) ? {srio_data[9:8],srio_data[39:11],3'b0} : {srio_data[23:0],10'b0};
  // Messaging fields
  assign msglen_bt1   = (DEVICEID_WIDTH == 8) ? srio_data[39:36] : srio_data[23:20];
  assign letter_bt1   = (DEVICEID_WIDTH == 8) ? srio_data[31:30] : srio_data[15:14];
  assign mbox_bt1     = (DEVICEID_WIDTH == 8) ? srio_data[29:28] : srio_data[13:12];
  assign msgseg_bt1   = (msglen_bt1 == 4'h0) ? 4'h0 : (DEVICEID_WIDTH == 8) ? srio_data[27:24] : srio_data[11:8];
  assign xmbox_bt1    = (msglen_bt1 != 4'h0) ? 4'h0 : (DEVICEID_WIDTH == 8) ? srio_data[27:24] : srio_data[11:8];

  // Extract the ssize for message transactions
  always @* begin
    case (sizestat_bt1)
      4'b1001: {bad_ssize,ssize_bt1} = 9'h0_07;
      4'b1010: {bad_ssize,ssize_bt1} = 9'h0_0F;
      4'b1011: {bad_ssize,ssize_bt1} = 9'h0_1F;
      4'b1100: {bad_ssize,ssize_bt1} = 9'h0_3F;
      4'b1101: {bad_ssize,ssize_bt1} = 9'h0_7F;
      4'b1110: {bad_ssize,ssize_bt1} = 9'h0_FF;
      default: {bad_ssize,ssize_bt1} = 9'h1_xx;
    endcase
  end

  // Create registered versions of header fields for transactions with >1 DWORD headers
  always @(posedge log_clk) begin
    // No reset needed because only sampled on valid data
    if (bufr_sof && bufr_active && !SHORT_HEADERS_ONLY) begin
      crf_bt2        <= #TCQ crf_bt1;
      prio_bt2       <= #TCQ prio_bt1;
      ttype_bt2      <= #TCQ ttype_bt1;
      rdwrsize_bt2   <= #TCQ sizestat_bt1;
      sizestat_bt2   <= #TCQ sizestat_bt1;
      tid_bt2        <= #TCQ tid_bt1;
      haddr_bt2      <= #TCQ haddr_bt1;
      ok_bt2         <= #TCQ ok_bt1;
      swr_haddr_bt2  <= #TCQ swr_addr_bt1[33:10];
    end
  end

  // Capture header fields always on the second DWORD
  assign swr_addr_bt2 = {srio_data[57:56],swr_haddr_bt2,srio_data[63:58],2'b0}; //Only needed for 16-bit device IDs
  assign laddr_bt2    = (DEVICEID_WIDTH == 8) ? srio_data[63:59] : srio_data[63:43];
  assign wdptr_bt2    = (DEVICEID_WIDTH == 8) ? srio_data[58]    : srio_data[42];
  assign xamsbs_bt2   = (DEVICEID_WIDTH == 8) ? srio_data[57:56] : srio_data[41:40];

  // Compute the HELLO size field and address lsbs for I/O transactions based on RapidIO Spec Part 1 Table 4-3/4
  // Note that some of the values below are not supported for writes but will not be flagged as "bad" (saves resources)
  always @* begin
    case({wdptr_bt2,rdwrsize_bt2})
      5'b1_0011: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h0_00; // 1 byte
      5'b1_0010: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h1_00; // 1 byte
      5'b1_0001: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h2_00; // 1 byte
      5'b1_0000: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h3_00; // 1 byte
      5'b0_0011: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h4_00; // 1 byte
      5'b0_0010: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h5_00; // 1 byte
      5'b0_0001: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h6_00; // 1 byte
      5'b0_0000: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h7_00; // 1 byte
      5'b1_0110: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h0_01; // 2 bytes
      5'b1_0100: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h2_01; // 2 bytes
      5'b0_0110: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h4_01; // 2 bytes
      5'b0_0100: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h6_01; // 2 bytes
      5'b1_0101: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h0_02; // 3 bytes
      5'b0_0101: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h5_02; // 3 bytes
      5'b1_1000: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h0_03; // 4 bytes
      5'b0_1000: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h4_03; // 4 bytes
      5'b1_0111: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h0_04; // 5 bytes
      5'b0_0111: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h3_04; // 5 bytes
      5'b1_1001: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h0_05; // 6 bytes
      5'b0_1001: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h2_05; // 6 bytes
      5'b1_1010: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h0_06; // 7 bytes
      5'b0_1010: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h1_06; // 7 bytes
      5'b0_1011: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h0_07; // 8 bytes
      5'b1_1011: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h0_0F; // 16 bytes
      5'b0_1100: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h0_1F; // 32 bytes
      5'b1_1100: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h0_3F; // 64 bytes
      5'b0_1101: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h0_5F; // 96 bytes - valid for reads only
      5'b1_1101: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h0_7F; // 128 bytes
      5'b0_1110: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h0_9F; // 160 bytes - valid for reads only
      5'b1_1110: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h0_BF; // 192 bytes - valid for reads only
      5'b0_1111: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h0_DF; // 224 bytes - valid for reads only
      5'b1_1111: {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'h0_FF; // 256 bytes
      default  : {bad_rdwrsize,addr_lsb_bt2,hello_size_bt2} = 12'b1_xxx_xxxxxxxx; // invalid size
    endcase
  end

  // Mask off size for maintenance responses
  assign maint_size_bt2 = (ftype_hold == FTYPE_MAINT[3:0]) && ttype_bt2[1] ? 8'b0 : hello_size_bt2;

  // Put the address together
  assign addr_bt2     = {xamsbs_bt2, haddr_bt2, laddr_bt2, addr_lsb_bt2};

  // Capture the FTYPE so that it's available after sof
  always @(posedge log_clk) begin
    // No reset needed because only sampled on valid data
    if (bufr_sof) begin
      ftype_hold     <= #TCQ ftype_bt1;
      ttype_hold     <= #TCQ ttype_bt1;
    end
  end

  // Create an FTYPE and a TTYPE bus that are valid throughout the packet
  assign bufr_ftype   = bufr_sof ? ftype_bt1 : ftype_hold;
  assign bufr_ttype   = bufr_sof ? ttype_bt1 : ttype_hold;

  // Create a flag to indicate whether the packet is being encoded into HELLO format
  always @* begin
    casex ({bufr_ftype,bufr_ttype})
      {FTYPE_NREAD,  4'b11xx}:  hello_encode = ENCODE_NREADATOMIC;
      {FTYPE_NREAD,  4'b0100}:  hello_encode = ENCODE_NREAD;
      {FTYPE_NWRITE, 4'b0100}:  hello_encode = ENCODE_NWRITE;
      {FTYPE_NWRITE, 4'b0101}:  hello_encode = ENCODE_NWRITE_R;
      {FTYPE_NWRITE, 4'b110x}:  hello_encode = ENCODE_NWRITEATOMIC;
      {FTYPE_NWRITE, 4'b1110}:  hello_encode = ENCODE_NWRITEATOMIC;
      {FTYPE_SWRITE, 4'bxxxx}:  hello_encode = ENCODE_SWRITE;
      {FTYPE_MAINT,  4'b00xx}:  hello_encode = ENCODE_MAINT;
      {FTYPE_DS,     4'bxxxx}:  hello_encode = ENCODE_DS;
      {FTYPE_DB,     4'bxxxx}:  hello_encode = ENCODE_DB;
      {FTYPE_MSG,    4'bxxxx}:  hello_encode = ENCODE_MSG;
      {FTYPE_RESP,   4'b0000}:  hello_encode = ENCODE_RESPNODATA;
      {FTYPE_RESP,   4'b1000}:  hello_encode = ENCODE_RESPWDATA;
      {FTYPE_RESP,   4'b0001}:  hello_encode = ENCODE_RESPMSG;
      default:                  hello_encode = 1'b0;
    endcase
  end

  // Register hello_encode to use after sof to ease timing
  always @(posedge log_clk) begin
    hello_encode_q <= #TCQ hello_encode;
  end

  // Mark the packet as an unsupported type if it's not enabled
  always @* begin
    casex ({bufr_ftype,bufr_ttype})
      {FTYPE_NREAD,  4'b11xx}:  unsupported_type_d = !TARGET_ATOMIC;
      {FTYPE_NREAD,  4'b0100}:  unsupported_type_d = !TARGET_NREAD;
      {FTYPE_NWRITE, 4'b0100}:  unsupported_type_d = !TARGET_NWRITE;
      {FTYPE_NWRITE, 4'b0101}:  unsupported_type_d = !TARGET_NWRITE_R;
      {FTYPE_NWRITE, 4'b110x}:  unsupported_type_d = !TARGET_ATOMIC;
      {FTYPE_NWRITE, 4'b1110}:  unsupported_type_d = !TARGET_ATOMIC;
      {FTYPE_SWRITE, 4'bxxxx}:  unsupported_type_d = !TARGET_SWRITE;
      {FTYPE_MAINT,  4'b00xx}:  unsupported_type_d = 1'b0;
      {FTYPE_DS,     4'bxxxx}:  unsupported_type_d = !TARGET_DS;
      {FTYPE_DB,     4'bxxxx}:  unsupported_type_d = !TARGET_DB;
      {FTYPE_MSG,    4'bxxxx}:  unsupported_type_d = !MSG_SINK_SINGLE && !MSG_SINK_MULTI;
      {FTYPE_RESP,   4'b0000}:  unsupported_type_d = !INIT_NWRITE_R   && !INIT_DB;
      {FTYPE_RESP,   4'b1000}:  unsupported_type_d = !INIT_NREAD      && !INIT_ATOMIC;
      {FTYPE_RESP,   4'b0001}:  unsupported_type_d = !MSG_INIT_SINGLE && !MSG_INIT_MULTI;
      default:                  unsupported_type_d = 1'b1;
    endcase
  end

  // }}} end Parse Received Packet


  // Short and Long header for ftype9
  
 reg [3:0] bufr_ftype_q;

  assign long_header_ftype9  = (FTYPE_DS == bufr_ftype_q) && (tid_bt2[7:6] != 2'b00) && (DEVICEID_WIDTH == 16);
  assign short_header_ftype9  = (FTYPE_DS == bufr_ftype) && (tid_bt1[7:6] == 2'b00) && (DEVICEID_WIDTH == 16);

  // {{{ Create HELLO Header and Data

generate if (DEVICEID_WIDTH == 8) begin: hello_rx_8devid_gen
  // Packets are different based on DEVICEID_WIDTH, so using a generate
  // in order to separate those cases
  always @* begin
    // On SOF:
    //  - Header is only valid if the header is <1 DWORD
    //  - Data is never valid
    if (bufr_sof) begin
      data_stage    = 1'b0;
      case (bufr_ftype)
        FTYPE_NREAD:    header_stage = 1'b0;
        FTYPE_NWRITE:   header_stage = 1'b0;
        FTYPE_SWRITE:   header_stage = 1'b1;
        FTYPE_MAINT:    header_stage = 1'b0;
        FTYPE_DS:       header_stage = 1'b1;
        FTYPE_MSG:      header_stage = 1'b1;
        FTYPE_DB:       header_stage = 1'b1;
        FTYPE_RESP:     header_stage = 1'b1;
        default:        header_stage = 1'b0;
      endcase

    // On the second beat:
    //  - Header is only valid if the header is >1 DWORD
    //  - Data is valid if header is not
    end else if (bufr_second) begin
      case (bufr_ftype)
        FTYPE_NREAD:    header_stage = 1'b1;
        FTYPE_NWRITE:   header_stage = 1'b1;
        FTYPE_SWRITE:   header_stage = 1'b0;
        FTYPE_MAINT:    header_stage = 1'b1;
        FTYPE_DS:       header_stage = 1'b0;
        FTYPE_MSG:      header_stage = 1'b0;
        FTYPE_RESP:     header_stage = 1'b0;
        default:        header_stage = 1'b0;
      endcase
      data_stage    =  !header_stage && hello_encode_q;

    // After the second beat:
    //  - Header is never valid
    //  - Data is always valid
    end else if (bufr_active && hello_encode_q) begin
      header_stage  = 1'b0;
      data_stage    = 1'b1;
    end else begin
      header_stage  = 1'b0;
      data_stage    = 1'b0;
    end
  end

  // Create the header
  always @* begin
    if (bufr_sof && !LONG_HEADERS_ONLY) begin
      case (bufr_ftype)
        FTYPE_NREAD:
          hello_header = 64'bx; // NREAD header will be valid on second beat
        FTYPE_NWRITE:
          hello_header = 64'bx; // NWRITE header will be valid on second beat
        FTYPE_SWRITE:
          hello_header = {8'b0,ftype_bt1,4'b0,1'b0,prio_bt1,crf_bt1,8'b0,1'b0,1'b0,swr_addr_bt1};
        FTYPE_MAINT:
          hello_header = 64'bx; // MAINT header will be valid on second beat
        FTYPE_DS:
          hello_header = {tid_bt1,ftype_bt1,4'b0,1'b0,prio_bt1,crf_bt1,ttype_bt1,sizestat_bt1,4'b0,haddr_bt1[23:8],haddr_bt1[23:8]};
        FTYPE_DB:
          hello_header = {tid_bt1,ftype_bt1,4'b0,1'b0,prio_bt1,crf_bt1,8'b0,1'b0,1'b0,2'b0,haddr_bt1[23:8],16'b0};
        FTYPE_MSG:
          hello_header = {msglen_bt1,msgseg_bt1,ftype_bt1,5'b0,prio_bt1,crf_bt1,ssize_bt1,1'b0,25'b0,xmbox_bt1,
                          mbox_bt1,2'b0,letter_bt1};
        FTYPE_RESP:
          hello_header = {tid_bt1,ftype_bt1,ttype_bt1,1'b0,prio_bt1,crf_bt1,8'b0,!ok_bt1,1'b0,2'b0,32'b0};
        default:
          hello_header = 64'bx;
      endcase
    end else if (!SHORT_HEADERS_ONLY) begin
      // NREAD, NWRITE, and MAINT all use the same header fields
      hello_header = {tid_bt2,ftype_hold,ttype_bt2,1'b0,prio_bt2,crf_bt2,maint_size_bt2,!ok_bt2,1'b0,addr_bt2};
    end else begin
      hello_header = 64'bx;
    end
  end

  // Create (shift) the data
  always @* begin
    case (bufr_ftype)
      FTYPE_NREAD:  begin
                	hello_data = {srio_data_hold[55:0],srio_data[63:56]};
			hello_tkeep = 8'hFF;
		      end
      FTYPE_NWRITE:  begin
		       	hello_data = {srio_data_hold[55:0],srio_data[63:56]};
			hello_tkeep = 8'hFF;
		      end
      FTYPE_SWRITE:   begin 
		      hello_data = {srio_data_hold[7:0], srio_data[63:8]};
			hello_tkeep = 8'hFF;
		      end
      FTYPE_MAINT:    begin 
		      hello_data = {srio_data_hold[55:0],srio_data[63:56]};
         		hello_tkeep = 8'hFF;
		      end

      FTYPE_DS:       begin 
                	hello_data = (tid_bt2[7:6] == 2'b00) ? {srio_data_hold[23:0],srio_data[63:24]} :
	                            {srio_data_hold[7:0],srio_data[63:8]};
                	hello_tkeep = (tid_bt2[7:6] == 2'b00) ? {srio_tkeep_hold[2:0],srio_tkeep[7:3]} :
	                            {srio_tkeep_hold[0],srio_tkeep[7:1]};
	        	end	  
	FTYPE_DB:       begin 
			hello_data = 64'bx; // There is never a data phase for DB transactions
         		hello_tkeep = 8'hFF;
		      end
     FTYPE_MSG:      begin 
		      hello_data = {srio_data_hold[23:0],srio_data[63:24]};
         		hello_tkeep = 8'hFF;
		      end
      FTYPE_RESP:     begin 
		      hello_data = {srio_data_hold[23:0],srio_data[63:24]};
         		hello_tkeep = 8'hFF;
		      end
      default:        begin 
		      hello_data = 64'bx;
         		hello_tkeep = 8'hFF;
		      end
    endcase
  end

end // end if (DEVICEID_WIDTH == 8)
// When using 16-bit device IDs, data alignment is different
else begin: hello_rx_16devid_gen // if (DEVICEID_WIDTH == 16)

  always @* begin
    // On SOF:
    //  - Header is only valid if the header is <1 DWORD
    //  - Data is never valid
    if (bufr_sof) begin
      case (bufr_ftype)
        FTYPE_NREAD:    header_stage = 1'b0;
        FTYPE_NWRITE:   header_stage = 1'b0;
        FTYPE_SWRITE:   header_stage = 1'b0;
        FTYPE_MAINT:    header_stage = 1'b0;
        FTYPE_DS:       header_stage = (tid_bt1[7:6] == 2'b00) ? 1'b1 : 1'b0;
        FTYPE_DB:       header_stage = 1'b0;
        FTYPE_MSG:      header_stage = 1'b1;
        FTYPE_RESP:     header_stage = 1'b1;
        default:        header_stage = 1'b0;
      endcase
      data_stage    = 1'b0;

    // On the second beat:
    //  - Header is only valid if the header is >1 DWORD
    //  - Data is valid if header is not
    end else if (bufr_second) begin
      case (bufr_ftype)
        FTYPE_NREAD:    header_stage = 1'b1;
        FTYPE_NWRITE:   header_stage = 1'b1;
        FTYPE_SWRITE:   header_stage = 1'b1;
        FTYPE_MAINT:    header_stage = 1'b1;
        FTYPE_DS:       header_stage = (tid_bt2[7:6] == 2'b00) ? 1'b0 : 1'b1;
        FTYPE_DB:       header_stage = 1'b1;
        FTYPE_MSG:      header_stage = 1'b0;
        FTYPE_RESP:     header_stage = 1'b0;
        default:        header_stage = 1'b0;
      endcase
      data_stage    = !header_stage && hello_encode_q;

    // After the second beat:
    //  - Header is never valid
    //  - Data is always valid
    end else if (bufr_active && hello_encode_q) begin
      header_stage  = 1'b0;
      data_stage    = 1'b1;
    end else begin
      header_stage  = 1'b0;
      data_stage    = 1'b0;
    end
  end

  // Create the header
  always @* begin
    if (bufr_sof && (!LONG_HEADERS_ONLY || short_header_ftype9)) begin
      case (bufr_ftype)
        FTYPE_NREAD:
          hello_header = 64'bx; // NREAD header not used on SOF
        FTYPE_NWRITE:
          hello_header = 64'bx; // NWRITE header not used on SOF
        FTYPE_SWRITE:
          hello_header = 64'bx; // SWRITE header not used on SOF
        FTYPE_MAINT:
          hello_header = 64'bx; // Maintenance header not used on SOF
        FTYPE_DS:
          hello_header = {tid_bt1,ftype_bt1,4'b0,1'b0,prio_bt1,crf_bt1,ttype_bt1,sizestat_bt1,4'b0,srio_data[23:8],srio_data[23:8]};
        FTYPE_DB:
          hello_header = 64'bx; // Doorbell header not used on SOF
        FTYPE_MSG:
          hello_header = {msglen_bt1,msgseg_bt1,ftype_bt1,5'b0,prio_bt1,crf_bt1,ssize_bt1,1'b0,25'b0,
                          xmbox_bt1,mbox_bt1,2'b0,letter_bt1};
        FTYPE_RESP:
          hello_header = {tid_bt1,ftype_bt1,ttype_bt1,1'b0,prio_bt1,crf_bt1,8'b0,!ok_bt1,1'b0,2'b0,32'b0};
        default:
          hello_header = 64'bx;
      endcase
    end else if (!SHORT_HEADERS_ONLY) begin
      case (bufr_ftype)
        FTYPE_NREAD:
          hello_header = {tid_bt2,ftype_hold,ttype_bt2,1'b0,prio_bt2,crf_bt2,hello_size_bt2,2'b0,addr_bt2};
        FTYPE_NWRITE:
          hello_header = {tid_bt2,ftype_hold,ttype_bt2,1'b0,prio_bt2,crf_bt2,hello_size_bt2,2'b0,addr_bt2};
        FTYPE_SWRITE:                                                                            //RSRV //XAMSBS                          
          hello_header = {8'b0,ftype_hold,4'b0,1'b0,prio_bt2,crf_bt2,8'b0,2'b0,swr_addr_bt2[33:3],1'b0,swr_addr_bt2[1:0]};
        FTYPE_MAINT:
          hello_header = {tid_bt2,ftype_hold,ttype_bt2,1'b0,prio_bt2,crf_bt2,maint_size_bt2,!ok_bt2,1'b0,addr_bt2};
        FTYPE_DS:
          hello_header = {tid_bt2,ftype_hold,4'b0,1'b0,prio_bt2,crf_bt2,ttype_bt2,sizestat_bt2,4'b0,haddr_bt2,srio_data[63:56],haddr_bt2,srio_data[63:56]};
        FTYPE_DB:
          hello_header = {tid_bt2,ftype_hold,4'b0,1'b0,prio_bt2,crf_bt2,8'b0,2'b0,2'b0,addr_bt2[31:16],16'b0};
        FTYPE_MSG:
          hello_header = 64'bx; // Message header only used on SOF
        FTYPE_RESP:
          hello_header = 64'bx; // Response header only used on SOF
        default:
          hello_header = 64'bx;
      endcase
    end else begin
      hello_header = 64'bx;
    end
  end

  // Create (shift) the data
  always @* begin
    case (bufr_ftype)

        FTYPE_NREAD:  begin
                        hello_data = {srio_data_hold[39:0],srio_data[63:40]};
			hello_tkeep = 8'hFF;
		      end
      FTYPE_NWRITE:  begin
                        hello_data = {srio_data_hold[39:0],srio_data[63:40]};
			hello_tkeep = 8'hFF;
		      end
      FTYPE_SWRITE:   begin 
                        hello_data = {srio_data_hold[55:0],srio_data[63:56]};
			hello_tkeep = 8'hFF;
		      end
      FTYPE_MAINT:    begin 
                        hello_data = {srio_data_hold[39:0],srio_data[63:40]};
         		hello_tkeep = 8'hFF;
		      end

      FTYPE_DS:       begin     
                	hello_data = (tid_bt2[7:6] == 2'b00) ? {srio_data_hold[7:0],srio_data[63:8]} :
	                            {srio_data_hold[55:0],srio_data[63:56]};
                	hello_tkeep = (tid_bt2[7:6] == 2'b00) ? {srio_tkeep_hold[0],srio_tkeep[7:1]} :
	                            {srio_tkeep_hold[6:0],srio_tkeep[7]};
			end
	FTYPE_DB:       begin 
			hello_data = 64'bx; // There is never a data phase for DB transactions
         		hello_tkeep = 8'hFF;
		      end
     FTYPE_MSG:      begin 
                        hello_data = {srio_data_hold[7:0],srio_data[63:8]};
         		hello_tkeep = 8'hFF;
		      end
      FTYPE_RESP:     begin 
                        hello_data = {srio_data_hold[7:0],srio_data[63:8]};
         		hello_tkeep = 8'hFF;
		      end
      default:        begin 
		      hello_data = 64'bx;
         		hello_tkeep = 8'hFF;
		      end

    endcase
  end

end endgenerate // end if (DEVICEID_WIDTH == 16)

  //*ASSERTION*
  //(ap_data_stage_x): data_stage should not be 1'bx when hello_encode is asserted
  //(ap_header_or_data_stage_for_hello): Either header_stage or data_stage is high during hello packet (except on sof)
  //(ap_not_header_and_data_stage): header_stage and data_stage do not assert simultaneously
  //(ap_hello_header_not_x): hello_header should not be x when header_stage is asserted
  //(ap_hello_data_not_x): hello_data should not be x when data_stage is asserted

  // }}} Create HELLO Header and Data

  // {{{ Output Generation
  // + {{{ Arbiter Interface +


  reg pkt_extend;
  wire pkt_end;
  reg bufr_active_q;


  assign pkt_extend_d = (pkt_extend && pkt_end) ? 1'b0 : (!arb_stall && hello_encode) ? ((long_header_ftype9 && bufr_last && srio_tkeep[6]) || (short_header_ftype9 && bufr_last && srio_tkeep[0])) : pkt_extend;
 
  assign pkt_end = pkt_extend && LE_lhrx_tvalid && LE_lhrx_tlast && LA_lhrx_tready; 



  always @(posedge log_clk) begin
    if (log_rst_q) begin
      pkt_extend <= #TCQ 1'b0;
      bufr_active_q <= #TCQ 1'b0;
      bufr_ftype_q <= #TCQ 4'b0000;
    end else begin
     pkt_extend <= pkt_extend_d;
     bufr_active_q <= bufr_active;
     bufr_ftype_q <= #TCQ bufr_ftype;
    end
  end



  // Create the tvalid signal
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LE_lhrx_tvalid <= #TCQ 1'b0;
    end else if (!arb_stall) begin
      if (!hello_encode && !pkt_extend) begin
        LE_lhrx_tvalid <= #TCQ bufr_active || (arb_stall_q && arb_stall_vld);
      end else begin
        LE_lhrx_tvalid <= #TCQ (bufr_active && (header_stage || data_stage)) || (arb_stall_q && arb_stall_vld && !pkt_end) || (pkt_extend && !pkt_end);
      end
    end
  end

  // Create the TDATA and TKEEP buses for the packet
  always @(posedge log_clk) begin
    if (!arb_stall) begin
      if (!hello_encode && !pkt_extend) begin
        LE_lhrx_tdata <= #TCQ bufr_data;
        LE_lhrx_tkeep <= #TCQ bufr_keep;
      end else if (header_stage && !pkt_extend) begin
        LE_lhrx_tdata <= #TCQ hello_header;
        LE_lhrx_tkeep <= #TCQ 8'hFF;
      end else if (data_stage || (arb_stall_q && !arb_stall_sof) || pkt_extend) begin
        LE_lhrx_tdata <= #TCQ pkt_extend  ? {srio_data_hold[55:0],8'h0} : hello_data;
        LE_lhrx_tkeep <= #TCQ pkt_extend ? {srio_tkeep_hold[6:0],1'b0} : hello_tkeep;

      end
    end
  end

  // Form the tuser bus for the packet, using the decoded src and dest IDs and the incoming tuser.
  // Register TUSER and the unsupported type indicator on SOF.
  always @(posedge log_clk) begin
    if (!arb_stall) begin
      if (bufr_sof) begin
        LE_lhrx_tuser       <= #TCQ {srcid_bt1,destid_bt1,bufr_user[7:6],hello_encode,bufr_user[4:0]};
      end
        LE_unsupported_type <= #TCQ unsupported_type_d && !(pkt_extend && !pkt_end);
    end
  end

  // Create the tlast signal for the packet
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LE_lhrx_tlast        <= #TCQ 1'b0;
    end else if (!arb_stall) begin
      LE_lhrx_tlast        <= #TCQ (bufr_last && (!hello_encode || header_stage || data_stage || arb_stall_q)
                                   && !pkt_extend_d) || (pkt_extend && !pkt_end) ;

    end
  end


  // Internal Coverage and Assertions
  //*COVERAGE*
  //(cp_lhrx_tlast_set_and_clr): The set and clear conditions for LE_lhrx_tlast happen together
  //(cp_lhrx_tvalid_set_and_clr): The set and clear conditions for LE_lhrx_tvalid happen together

  // Arbiter Interface Coverage and Assertions
  //*COVERAGE*
  //(cp_lhrx_b2b_single_cycle): There are back-to-back single-cycle packets on the lhrx interface

  //*ASSERTION*
  //(ap_lhrx_valid_high_until_active): Once asserted, LE_lhrx_tvalid stays high until LA_lhrx_tready is asserted
  //(ap_no_x_on_lhrx_tvalid): When LE_lhrx_tvalid is asserted, other outputs cannot be unknown

  // + }}} end Arbiter Interface +

  // + {{{ Buffer Interface +

  // Use the arbiter's ready signal as the bufr_ready to avoid adding a lot of shadow registers
 
  assign LE_bufr_tready = LA_lhrx_tready && !((bufr_ftype == 4'h9) && bufr_last && !bufr_last_q) && !pkt_extend_d;

  // RX Buffer Interface Coverage and Assertions
  //*COVERAGE*
  //(cp_bufr_valid_drops_mid_packet): The receive buffer stalls mid-packet
  //(cp_bufr_valid_drops_after_sof): The receive buffer stalls on the second beat
  //(cp_bufr_valid_drops_between_packets): The receive buffer stalls between packets
  //(cp_bufr_ready_drops_mid_packet): The hello_encoder stalls mid-packet
  //(cp_bufr_ready_drops_after_sof): The hello_encoder stalls on the second beat
  //(cp_bufr_ready_drops_between_packets): The hello_encoder stalls between packets
  //(cp_rx_b2b_two_single_cycle_pkts): cover that back to back single cycle packets exit the buffer

  //*ASSERTION*
  //(ap_bufr_valid_high_until_active): Once asserted, BR_bufr_tvalid stays high until LE_bufr_tready is asserted
  //(ap_bufr_keep_ff_w_valid): for every valid cycle other that last the strobe must be 'FF

  // + }}} end Buffer Interface +
  // }}} Output Generation

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/log/log_hello/srio_gen2_v4_1_16_hello_decoder.v#4 $
//----------------------------------------------------------------------
//
// HELLO_DECODER
// Description:
// This module converts packets from HELLO format and sRIO Native format
// to Buffer Native format. It sits in the LOG TX data path between the
// LOG TX Arbiter and the TX Buffer
//
// Hierarchy:
// LOG_TOP
//    |___HELLO_DECODER - this module
// ---------------------------------------------------------------------

`timescale 1ps/1ps

// ------------------------------------------------
// below attribute is added to supress the synthesis warnings in vivado tool 8:3332
(* DowngradeIPIdentifiedWarnings="yes" *)
// ------------------------------------------------

module srio_gen2_v4_1_16_hello_decoder
#(
  parameter TCQ            =  100, // in ps
  parameter DEVICEID_WIDTH =    8, // Indicates Source/Dest ID width {8, 16}
  parameter DECODE_FT02    =    1, // If 1, must be able to decode FTYPE2 (NREAD and ATOMIC) {0, 1}
  parameter DECODE_FT05    =    1, // If 1, must be able to decode FTYPE5 (NWRITE, NWRITE_R, and ATOMIC) {0, 1}
  parameter DECODE_FT06    =    1, // If 1, must be able to decode FTYPE6 (SWRITE) {0, 1}
  parameter DECODE_FT08    =    1, // If 1, must be able to decode FTYPE8 (MAINTENANCE) {0, 1}
  parameter DECODE_FT09    =    1, // If 1, must be able to decode FTYPE9 (DATA STREAMING) {0, 1}
  parameter DECODE_FT10    =    1, // If 1, must be able to decode FTYPE10 (DOORBELL) {0, 1}
  parameter DECODE_FT11    =    1, // If 1, must be able to decode FTYPE11 (MESSAGE) {0, 1}
  parameter DECODE_FT13    =    1, // If 1, must be able to decode FTYPE13 (RESPONSE) {0, 1}  
  parameter CRF_SUPPORT    =    1) // The CRF support parameter set from the GUI top // CR# 820838
(
  // {{{ Port Declarations
  // System Signals
  input                         log_clk,
  input                         log_rst,

  // TX Buffer Interface
  output reg                    LD_buft_tvalid,       // Valid Packet Beat
  input                         BT_buft_tready,       // Packet Beat Accepted
  output reg [63:0]             LD_buft_tdata = 0,    // Packet Data
  output reg [7:0]              LD_buft_tkeep = 0,    // Valid bytes in this beat, only valid on last
  output reg                    LD_buft_tlast = 0,    // Last Beat
  output reg [7:0]              LD_buft_tuser = 0,    // {DEST_ID, SRC_ID, 3'h0, RESPONSE, 1'b0, VC, CRF, 1'b0}

  // LOG Arbiter Interface
  input                         LA_lhtx_tvalid,       // Valid Packet Beat
  output reg                    LD_lhtx_tready = 0,   // Packet Beat Accepted
  input      [63:0]             LA_lhtx_tdata,        // Packet Data
  input      [7:0]              LA_lhtx_tkeep,        // Valid bytes in this beat, only valid on last
  input                         LA_lhtx_tlast,        // Last Beat
  input      [39:0]             LA_lhtx_tuser         // {DEST_ID, SRC_ID, 2'h0, HELLO_FMT, RESPONSE, 1'b0, VC, CRF, 1'b0}

  // }}} end Port Declarations
);

 // {{{ Local Parameters
  // Spec defined parameters
  // ------------------------------------------------------------
  // Ftype (plus 16 if not supported - used in packet decode case statements)
  localparam [4:0] FTYPE_NREAD      = {(DECODE_FT02 == 0),4'b0010};
  localparam [4:0] FTYPE_NWRITE     = {(DECODE_FT05 == 0),4'b0101};
  localparam [4:0] FTYPE_SWRITE     = {(DECODE_FT06 == 0),4'b0110};
  localparam [4:0] FTYPE_MAINT      = {(DECODE_FT08 == 0),4'b1000};
  localparam [4:0] FTYPE_DS         = {(DECODE_FT09 == 0),4'b1001};
  localparam [4:0] FTYPE_DB         = {(DECODE_FT10 == 0),4'b1010};
  localparam [4:0] FTYPE_MSG        = {(DECODE_FT11 == 0),4'b1011};
  localparam [4:0] FTYPE_RESP       = {(DECODE_FT13 == 0),4'b1101};
  localparam [4:0] TTYPE_MSGRESP    = {(DECODE_FT11 == 0),4'b0001};
  // tt field for outgoing packets (spec Rev 2.1 Part 3 Section 2.4)
  localparam TT                     = (DEVICEID_WIDTH == 8) ? 2'b0 : 2'b01;
  // }}} end Local Parameters

  // {{{ Wire Declarations
  reg           log_rst_q = 1;

  wire          lhtx_active;        // Transfer on lhtx (TVALID and TREADY asserted)
  reg           lhtx_tlast_hold = 1;// The lhtx_tlast input captured on lhtx_active for creating sof signal
  reg [7:0]     lhtx_tkeep_hold = 1;// The lhtx_tlast input captured on lhtx_active for creating sof signal
  reg           lhtx_sof_hold;      // The sof signal captured on lhtx_active for creating the second beat indicator
  wire          lhtx_sof;           // The start-of-frame on the lhtx interface is transferred
  wire          lhtx_second;        // The second beat on the lhtx interface is transferred
  reg           hello_fmt;          // The packet received from the arbiter is in HELLO format
  wire          hello_decode;       // The current packet will be decoded from HELLO
  wire [15:0]   hello_srcid;        // The Source ID from the TUSER input
  wire [15:0]   hello_destid;       // The Destination ID from the TUSER input
  wire [7:0]    hello_tid;          // The TID for the HELLO packet
  wire [3:0]    hello_ftype;        // The FTYPE for the HELLO packet
  wire [3:0]    hello_ttype;        // The TTYPE for the HELLO packet
  wire          hello_vc;           // The VC bit for the HELLO packet
  wire [1:0]    hello_prio;         // The priority field for the HELLO packet
  wire          hello_crf;          // The CRF bit for the HELLO packet
  wire [7:0]    hello_size;         // The size of the packet in HELLO format (Number of bytes minus 1)
  wire [3:0]    hello_stat;         // The HELLO status expanded into sRIO format (4'b0000 - OK/DONE, 4'b0111 - ERR)
  wire [1:0]    hello_xamsbs;       // The xamsbs field derived from the address and size fields
  wire [31:0]   hello_addr;         // The address (or config offset) for the HELLO packet, minus the xamsbs
  wire          hello_maintresp;    // The HELLO packet is a maint response
  reg           bad_rdwrsize;       // The rdsize/wrsize decode detected an invalid addr/size combo
  reg           hello_wdptr;        // The wdptr value for the packet after conversion to sRIO Native
  reg  [3:0]    hello_rdwrsize;     // The rdsize or wrsize value decoded from the address and size
  wire [3:0]    hello_sizestat;     // The size/status field used for
  reg           bad_ssize;          // Unable to decode a valid ssize for a message transaction
  reg  [3:0]    hello_ssize;        // The ssize for a message transaction
  wire [3:0]    hello_msglen;       // The msglen field for a message
  wire [1:0]    hello_letter;       // The letter field for a message
  wire [1:0]    hello_mbox;         // The mbox field for a message
  wire [3:0]    hello_msgseg;       // The msgseg field for a message
  wire [3:0]    hello_xmbox;        // The xmbox field for a message
  wire [3:0]    hello_msgsegxmbox;  // A mux of the msgseg and xmbox based on msg length
  reg  [1:0]    hello_xamsbs_hold;  // hello_xamsbs captured on lhtx_active for use in the second DWORD
  reg  [23:0]   hello_addr_hold;    // hello_addr captured on lhtx_active for use in the second DWORD
  reg  [63:0]   hello_data_hold;    // LA_lhtx_tdata captured on lhtx_active for use in the subsequent DWORD
  reg           hello_wdptr_hold;   // hello_wdptr captured on lhtx_active for use in the second DWORD
  reg  [3:0]    lhtx_ftype_hold = 0;// hello_ftype captured on lhtx_sof so that it's available throughout the packet
  wire [3:0]    lhtx_ftype;         // FTYPE, valid throughout packet including sof
  wire          need_extra_beat;    // A beat needs to be inserted if the packet is more cycles on buft than lhtx
  reg           hd_insert_beat;     // Register extra beat request and hold through a stall (if applicable)
  wire          hd_insert_beat_clr; // The extra beat has been inserted
  wire          hd_update;          // The decoded data should be updated on the buft interface only if valid
  (* max_fanout = 50 *)             // added to meet the timings, 25/2/2015
  reg           hd_first = 1;       // Create a first beat indicator that is registered for the decoder
  (* max_fanout = 50 *)             // added to meet the timings, 25/2/2015
  reg           hd_second = 0;      // Create a second beat indicator that is registered for the decoder
  reg  [7:0]    hd_keep;            // The HELLO decoded keep signal which will be used to form TKEEP to the buffer
  reg  [63:0]   hd_data;            // The HELLO decoded data signal which will be used to form TDATA to the buffer
  reg  [7:0]    hd_user;            // The HELLO decoded user signal which will be used to form TUSER to the buffer
  reg           hd_last;            // The HELLO decoded last signal which will be used to form TLAST to the buffer
  reg  [7:0]    hd_we;              // A byte-wise write enable for the data bus for the output register
  reg           hd_vld;             // An indicator that the TVALID for the corresponding hd_data should be asserted
  wire [3:0]    srio_ftype;         // FTYPE of incoming sRIO Native packet (valid on lhtx_sof)
  wire [3:0]    srio_ttype;         // TTYPE of incoming sRIO Native packet (valid on lhtx_sof)
  wire          srio_resp;          // Decode sRIO Native pkt type to set RESPONSE bit in TUSER
  wire [7:0]    bn_keep;            // keep signal for decoded packet after Buffer Native conversion
  wire [63:0]   bn_data;            // data signal for decoded packet after Buffer Native conversion
  wire [7:0]    bn_we;              // Buffer Native byte-wise write en for the output data for HELLO decoded pkt
  wire [7:0]    buft_keep;          // keep signal after Buffer Native conversion or incoming keep if un-decoded type
  wire [63:0]   buft_data;          // data signal after Buffer Native conversion or incoming data if un-decoded type
  wire [7:0]    buft_user;          // user signal after Buffer Native conversion or incoming user if un-decoded type
  wire          buft_last;          // last signal after Buffer Native conversion or incoming last if un-decoded type
  wire [7:0]    buft_we;            // Byte-wise write en for the output data after muxing input and decoded stream
  wire          buft_vld;           // Valid indicator after muxing decoded pkt and input stream based on hello_decode
  wire          buffer_stall;       // The buffer is stalling the transmit data
  reg           buffer_stall_q;     // A registered version of buffer_stall used to find the falling edge
  wire          buffer_stall_fell;  // The falling edge of buffer_stall
  reg           buffer_stall_fell_q;// A registered version of buffer_stall_fell used for inserted beat after stall
  reg           buffer_stall_active;// The lhtx interface was active on the rising edge of buffer_stall
  reg           buffer_stall_valid; // The data was valid on the rising edge of buffer_stall
  reg           buffer_stall_sof;   // The data was an sof on the rising edge of buffer_stall
  reg           buffer_stall_last;  // The data for the buffer was the last beat on the rising edge of buffer_stall
  reg  [7:0]    holdreg_tkeep = 0;  // A shadow register for TKEEP for a buffer stall to preserve 1 cycle latency
  reg  [7:0]    holdreg_tuser = 0;  // A shadow register for TUSER for a buffer stall to preserve 1 cycle latency
  reg  [63:0]   holdreg_tdata = 0;  // A shadow register for TDATA for a buffer stall to preserve 1 cycle latency
  wire          ld_buft_tlast_d;    // Form TLAST for buft interface
  wire          ld_buft_tvalid_d;   // Form TVALID for buft interface
  // }}} end Wire Declarations


  // {{{ Register Reset
  // Must register the reset before use to reduce fanout
  always @(posedge log_clk) begin
    log_rst_q <= #TCQ log_rst;
  end
  // }}} end Register Reset

  // {{{ Create Control Signals

  // Track when data is transferred from the arbiter
  assign lhtx_active = LA_lhtx_tvalid && LD_lhtx_tready;

  // Keep track of first beat of data
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lhtx_tlast_hold <= #TCQ 1'b1; // Reset to one so that sof asserts for the first frame
      lhtx_sof_hold   <= #TCQ 1'b0;
      lhtx_tkeep_hold <= #TCQ 8'b1111_1111;
    end else if (lhtx_active) begin
      lhtx_tlast_hold <= #TCQ LA_lhtx_tlast;
      lhtx_sof_hold   <= #TCQ lhtx_sof;
      lhtx_tkeep_hold <= #TCQ LA_lhtx_tkeep;
    end
  end

  // Create sof indicator for lhtx interface
  assign lhtx_sof    = lhtx_active && lhtx_tlast_hold;

  // Create second beat indicator
  assign lhtx_second = ((lhtx_active && !lhtx_tlast_hold) || hd_insert_beat) && lhtx_sof_hold;

  // The packet is in HELLO format if bit 5 of the user field is set
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      hello_fmt <= #TCQ 1'b0;
    end else if (lhtx_sof) begin
      hello_fmt <= #TCQ LA_lhtx_tuser[5];
    end
  end

  // Indicate whether the packet is in HELLO format, valid throughout the packet (including on sof)
  assign hello_decode = lhtx_sof ? LA_lhtx_tuser[5] : hello_fmt;

  // Indicate when the Buffer is not accepting the data from the hello_decoder
  assign buffer_stall = LD_buft_tvalid && !BT_buft_tready;

  // Register buffer_stall flag so that falling edge can be detected
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      buffer_stall_q <= #TCQ 1'b0;
    end else begin
      buffer_stall_q <= #TCQ buffer_stall;
    end
  end

  // Indicate that the Buffer released the stall condition
  assign buffer_stall_fell = buffer_stall_q && !buffer_stall;

  // Register buffer_stall_fell flag for the special case where the buf stalls on the cycle before a beat is inserted
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      buffer_stall_fell_q <= #TCQ 1'b0;
    end else begin
      buffer_stall_fell_q <= #TCQ buffer_stall_fell;
    end
  end

  // Capture the state of the lhtx interface on a buffer stall to act accordingly when the stall releases
  // Need separate buffer_stall active and valid indicators because of MSGs and SWRITEs, which may not be vld on sof
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      buffer_stall_valid  <= #TCQ 1'b0;
      buffer_stall_active <= #TCQ 1'b0;
      buffer_stall_sof    <= #TCQ 1'b0;
      buffer_stall_last   <= #TCQ 1'b0;
    end else if (buffer_stall && !buffer_stall_q) begin
      buffer_stall_valid  <= #TCQ buft_vld && (lhtx_active || hd_insert_beat);
      buffer_stall_active <= #TCQ lhtx_active;
      buffer_stall_sof    <= #TCQ lhtx_sof;
      buffer_stall_last   <= #TCQ buft_last && (lhtx_active || hd_insert_beat);
    end
  end

  // }}} end Create Control Signals

  // {{{ Parse HELLO Packet

  // Extract header fields from TUSER bus on the arbiter interface
  assign hello_srcid     = LA_lhtx_tuser[39:24];
  assign hello_destid    = LA_lhtx_tuser[23:8];

  // Extract header fields from the TDATA bus on the arbiter interface
  assign hello_tid       = LA_lhtx_tdata[63:56];
  assign hello_ftype     = LA_lhtx_tdata[55:52];
  assign hello_ttype     = LA_lhtx_tdata[51:48];
  //FIXVC - VC bit is TBD - tdata[47]?
  assign hello_vc        = 1'b0;
  assign hello_prio      = LA_lhtx_tdata[46:45];

  generate if (CRF_SUPPORT == 1) // CR# 820838 
  begin: crf_included_decoder_gen
  assign hello_crf       = LA_lhtx_tdata[44];
  end 
  endgenerate

  generate if (CRF_SUPPORT == 0) // CR# 820838
  begin: crf_excluded_decoder_gen
      assign hello_crf       = 1'b0;
  end 
  endgenerate
  
  assign hello_size      = LA_lhtx_tdata[43:36];
  assign hello_stat      = {1'b0, {3{LA_lhtx_tdata[35]}} };
  assign hello_xamsbs    = LA_lhtx_tdata[33:32];
  assign hello_addr      = LA_lhtx_tdata[31:0];
  assign hello_maintresp = ({1'b0,hello_ftype} == FTYPE_MAINT) && (hello_ttype[3:1] == 3'b001);

  // Compute the RDSIZE/WRSIZE fields for I/O transactions based on RapidIO Spec Part 1 Table 4-3/4
  // Note that some of the values below are not supported for writes but will not be flagged as "bad" (saves resources)
  // "bad_rdwrsize" is informational for debug and is not used to create an error
  always @* begin
    case ({hello_addr[2:0],hello_size})
      11'h0_00: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_1_0011;
      11'h1_00: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_1_0010;
      11'h2_00: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_1_0001;
      11'h3_00: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_1_0000;
      11'h4_00: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_0_0011;
      11'h5_00: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_0_0010;
      11'h6_00: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_0_0001;
      11'h7_00: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_0_0000;
      11'h0_01: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_1_0110;
      11'h2_01: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_1_0100;
      11'h4_01: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_0_0110;
      11'h6_01: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_0_0100;
      11'h0_02: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_1_0101;
      11'h5_02: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_0_0101;
      11'h0_03: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_1_1000;
      11'h4_03: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_0_1000;
      11'h0_04: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_1_0111;
      11'h3_04: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_0_0111;
      11'h0_05: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_1_1001;
      11'h2_05: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_0_1001;
      11'h0_06: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_1_1010;
      11'h1_06: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_0_1010;
      11'h0_07: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_0_1011;
      11'h0_0F: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_1_1011;
      11'h0_1F: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_0_1100;
      11'h0_3F: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_1_1100;
      11'h0_5F: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_0_1101; // Valid for reads only
      11'h0_7F: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_1_1101;
      11'h0_9F: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_0_1110; // Valid for reads only
      11'h0_BF: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_1_1110; // Valid for reads only
      11'h0_DF: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_0_1111; // Valid for reads only
      11'h0_FF: {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b0_1_1111;
      default : {bad_rdwrsize,hello_wdptr,hello_rdwrsize} = 6'b1_0_0000;
    endcase
  end

  //*ASSERTION*
  //(ap_lhtx_valid_size_addr): Should only get valid size/address combos for MAINT reqs, NREADs and NWRITEs

  // Mux between size and status based on packet type (status for mant response, else size)
  assign hello_sizestat = hello_maintresp ? hello_stat : hello_rdwrsize;

  // Compute the SSIZE field for message transactions
  // "bad_ssize" is informational for debug and is not used to create an error
  always @* begin
    case (hello_size)
      8'h07  : {bad_ssize,hello_ssize} = 5'b0_1001;
      8'h0F  : {bad_ssize,hello_ssize} = 5'b0_1010;
      8'h1F  : {bad_ssize,hello_ssize} = 5'b0_1011;
      8'h3F  : {bad_ssize,hello_ssize} = 5'b0_1100;
      8'h7F  : {bad_ssize,hello_ssize} = 5'b0_1101;
      8'hFF  : {bad_ssize,hello_ssize} = 5'b0_1110;
      default: {bad_ssize,hello_ssize} = 5'b1_0000;
    endcase
  end

  //*ASSERTION*
  //(ap_lhtx_valid_ssize): Should only get valid size/address combos for Messages

  // Create the messaging fields in sRIO Native format
  assign hello_msglen      = LA_lhtx_tdata[63:60];
  assign hello_msgseg      = LA_lhtx_tdata[59:56];
  assign hello_xmbox       = LA_lhtx_tdata[9:6];
  assign hello_mbox        = LA_lhtx_tdata[5:4];
  assign hello_letter      = LA_lhtx_tdata[1:0];
  assign hello_msgsegxmbox = (hello_msglen == 4'h0) ? hello_xmbox : hello_msgseg;

  // Register header fields needed for the second DWORD
  always @(posedge log_clk) begin
   if (lhtx_active) begin
      hello_xamsbs_hold   <= #TCQ hello_xamsbs;
      hello_addr_hold     <= #TCQ (hello_maintresp == 1'b0) ? hello_addr[23:0] : 24'b0;
      hello_data_hold     <= #TCQ LA_lhtx_tdata;
      hello_wdptr_hold    <= #TCQ hello_wdptr;
    end
  end

  reg [7:0] lhtx_tid_hold;
  // Capture the FTYPE so that it's available after sof
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lhtx_ftype_hold     <= #TCQ 4'b0;
      lhtx_tid_hold     <= #TCQ 8'b0;
    end else if (lhtx_sof) begin
      lhtx_ftype_hold     <= #TCQ hello_ftype;
      lhtx_tid_hold     <= #TCQ hello_tid;
    end else if (ld_buft_tlast_d && !buffer_stall_q) begin
      lhtx_ftype_hold     <= #TCQ 4'b0;
      lhtx_tid_hold     <= #TCQ 8'b0;
    end
  end

  // Create a signal that will indicate the packet's FTYPE throughout the transfer on LHTX
  assign lhtx_ftype = (hd_first == 1) ? hello_ftype : lhtx_ftype_hold; // In (hd_first == 1) sttement, replaced case equality operator (===) with the logical equality (==) operator. CR 725563 fixed.
 
  // }}} end Parse HELLO Packet

  // {{{ Create sRIO Native packet
  // Build the sRIO Native packet from the HELLO packet

  // A beat needs to be inserted if the packet is longer on the buft interface than the lhtx
  assign need_extra_beat = LA_lhtx_tlast && lhtx_active && !buft_last;

  // Clear the insert beat request 
  assign hd_insert_beat_clr = !buffer_stall && (!buffer_stall_fell || buffer_stall_last);
  
  // Register the extra beat request, clearing after a stall (if applicable)
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      hd_insert_beat     <= #TCQ 1'b0;
    end else if (need_extra_beat) begin
      hd_insert_beat     <= #TCQ 1'b1;
    end else if (hd_insert_beat_clr) begin
      hd_insert_beat     <= #TCQ 1'b0;
    end
  end

  // Only update the data if the new data is fresh or an extra beat is needed to finish the packet
  assign hd_update = hd_insert_beat || lhtx_active;

  // Create a speculative sof indicator to ease timing of HELLO decode
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      hd_first     <= #TCQ 1'b1; // Reset to one so that hd_first is asserted for first packet
    end else if (LA_lhtx_tlast && lhtx_active && buft_last) begin // no extra beat needed for this packet - last=last
      hd_first     <= #TCQ 1'b1;
    end else if (hd_insert_beat && hd_insert_beat_clr) begin //insert_beat falling
      hd_first     <= #TCQ 1'b1;
    end else if (lhtx_active) begin
      hd_first     <= #TCQ 1'b0;
    end
  end

  // Create a speculative second beat indicator to ease timing of HELLO decode
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      hd_second     <= #TCQ 1'b0;
    end else if (lhtx_active && lhtx_sof && (!LA_lhtx_tlast || need_extra_beat)) begin
      hd_second     <= #TCQ 1'b1;
    end else if (lhtx_active || (hd_insert_beat && hd_insert_beat_clr)) begin
      hd_second     <= #TCQ 1'b0;
    end
  end

generate if (DEVICEID_WIDTH == 8) begin: hello_decoder_8devid_gen
  // Packets are different based on DEVICEID_WIDTH, so using a generate
  // in order to separate those cases
  always @* begin
    case ({1'b0,lhtx_ftype})
      FTYPE_NREAD,FTYPE_NWRITE: begin
        case ({hd_first,hd_second})
          2'b10: begin
            hd_keep = 8'b1111_1111;
            hd_data = {hello_prio,TT,hello_ftype,hello_destid[7:0],hello_srcid[7:0],hello_ttype,
                       hello_rdwrsize,hello_tid,hello_addr[31:8]};
            hd_user = {3'b0,1'b0,1'b0,hello_vc,hello_crf,1'b0};
            hd_last = 1'b0;
            hd_we   = 8'b1111_1111;
            hd_vld  = 1'b1;
          end
          2'b01: begin
            hd_keep = lhtx_tlast_hold ? 8'b1000_0000 : 8'b1111_1111;
            hd_data = {hello_addr_hold[7:3],hello_wdptr_hold,hello_xamsbs_hold,LA_lhtx_tdata[63:8]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = lhtx_tlast_hold;
            hd_we   = 8'b1111_1111;
            hd_vld  = 1'b1;
          end
          default: begin
            hd_keep = lhtx_tlast_hold ? 8'b1000_0000 : 8'b1111_1111;
            hd_data = {hello_data_hold[7:0],LA_lhtx_tdata[63:8]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = lhtx_tlast_hold;
            hd_we   = hd_update ? 8'b1111_1111 : 8'b0000_0000;
            hd_vld  = hd_update;
          end
        endcase
      end
      FTYPE_SWRITE: begin
        case ({hd_first,hd_second})
          2'b10: begin
            hd_keep = 8'b1111_1111;
            hd_data = {hello_prio,TT,hello_ftype,hello_destid[7:0],hello_srcid[7:0],
                       hello_addr[31:3],1'b0,hello_xamsbs, 8'bx};
            hd_user = {3'b0,1'b0,1'b0,hello_vc,hello_crf,1'b0};
            hd_last = 1'b0;
            hd_we   = 8'b1111_1110;
            hd_vld  = 1'b0;
          end
          2'b01: begin
            hd_keep = 8'b1111_1111;
            hd_data = {56'bx,LA_lhtx_tdata[63:56]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = 1'b0;
            hd_we   = 8'b0000_0001;
            hd_vld  = 1'b1;
          end
          default: begin
            hd_keep = lhtx_tlast_hold ? 8'b1111_1110 : 8'b1111_1111;
            hd_data = {hello_data_hold[55:0],LA_lhtx_tdata[63:56]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = lhtx_tlast_hold;
            hd_we   = hd_update ? 8'b1111_1111 : 8'b0000_0000;
            hd_vld  = hd_update;
          end
        endcase
      end
      FTYPE_MAINT: begin
        case ({hd_first,hd_second})
          2'b10: begin
            hd_keep = 8'b1111_1111;
            hd_data = {hello_prio,TT,hello_ftype,hello_destid[7:0],hello_srcid[7:0],hello_ttype,
                       hello_sizestat,hello_tid,hello_addr[31:8]};
            hd_user = {3'b0,hello_maintresp,1'b0,hello_vc,hello_crf,1'b0};
            hd_last = 1'b0;
            hd_we   = 8'b1111_1111;
            hd_vld  = 1'b1;
          end
          2'b01: begin
            hd_keep = lhtx_tlast_hold ? 8'b1000_0000 : 8'b1111_1111;
            hd_data = {hello_addr_hold[7:3],hello_wdptr_hold,2'b0,LA_lhtx_tdata[63:8]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = lhtx_tlast_hold;
            hd_we   = 8'b1111_1111;
            hd_vld  = 1'b1;
          end
          default: begin
            hd_keep = lhtx_tlast_hold ? 8'b1000_0000 : 8'b1111_1111;
            hd_data = {hello_data_hold[7:0],LA_lhtx_tdata[63:8]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = lhtx_tlast_hold;
            hd_we   = hd_update ? 8'b1111_1111 : 8'b0000_0000;
            hd_vld  = hd_update;
          end
        endcase
      end
      FTYPE_MSG: begin
        case ({hd_first,hd_second})
          2'b10: begin
            hd_keep = 8'b1111_1111;
            hd_data = {hello_prio,TT,hello_ftype,hello_destid[7:0],hello_srcid[7:0],hello_msglen,
                       hello_ssize,hello_letter,hello_mbox,hello_msgsegxmbox,24'bx};
            hd_user = {3'b0,1'b0,1'b0,hello_vc,hello_crf,1'b0};
            hd_last = 1'b0;
            hd_we   = 8'b1111_1000;
            hd_vld  = 1'b0;
          end
          2'b01: begin
            hd_keep = 8'b1111_1111;
            hd_data = {40'bx,LA_lhtx_tdata[63:40]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = 1'b0;
            hd_we   = 8'b0000_0111;
            hd_vld  = 1'b1;
          end
          default: begin
            hd_keep = lhtx_tlast_hold ? 8'b1111_1000 : 8'b1111_1111;
            hd_data = {hello_data_hold[39:0],LA_lhtx_tdata[63:40]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = lhtx_tlast_hold;
            hd_we   = hd_update ? 8'b1111_1111 : 8'b0000_0000;
            hd_vld  = hd_update;
          end
        endcase
      end
      FTYPE_DB: begin
            hd_keep = 8'b1111_1110;
            hd_data = {hello_prio,TT,hello_ftype,hello_destid[7:0],hello_srcid[7:0],
                       8'b0,hello_tid,hello_addr[31:16],8'bx};
            hd_user = {3'b0,1'b0,1'b0,hello_vc,hello_crf,1'b0};
            hd_last = 1'b1;
            hd_we   = 8'b1111_1110;
            hd_vld  = hd_update;
      end
      FTYPE_RESP: begin
        case ({hd_first,hd_second})
          2'b10: begin
            hd_keep = LA_lhtx_tlast ? 8'b1111_1000 : 8'b1111_1111;
            hd_data = {hello_prio,TT,hello_ftype,hello_destid[7:0],hello_srcid[7:0],hello_ttype,hello_stat,
                       hello_tid,24'bx};
            hd_user = {3'b0,1'b1,1'b0,hello_vc,hello_crf,1'b0};
            hd_last = LA_lhtx_tlast;
            hd_we   = 8'b1111_1000;
            hd_vld  = LA_lhtx_tlast;
          end
          2'b01: begin
            hd_keep = 8'b1111_1111;
            hd_data = {40'bx,LA_lhtx_tdata[63:40]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = 1'b0;
            hd_we   = 8'b0000_0111;
            hd_vld  = 1'b1;
          end
          default: begin
            hd_keep = lhtx_tlast_hold ? 8'b1111_1000 : 8'b1111_1111;
            hd_data = {hello_data_hold[39:0],LA_lhtx_tdata[63:40]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = lhtx_tlast_hold;
            hd_we   = hd_update ? 8'b1111_1111 : 8'b0000_0000;
            hd_vld  = hd_update;
          end
        endcase
      end
      FTYPE_DS: begin
        case ({hd_first,hd_second})
          2'b10: begin
            hd_keep = 8'b1111_1111;
            hd_data = {hello_prio,TT,hello_ftype,hello_destid[7:0],hello_srcid[7:0],hello_size,
                       hello_tid,(hello_tid[7:6] == 2'b01 ? hello_addr[15:0] : hello_addr[31:16]),8'bx};
            hd_user = {3'b0,1'b0,1'b0,hello_vc,hello_crf,1'b0};
            hd_last = 1'b0;
            hd_we   = (hello_tid[7:6] == 2'b00) ? 8'b1111_1000 : 8'b1111_1110;
            hd_vld  = 1'b0;
          end
          2'b01: begin
            hd_keep = 8'b1111_1111;
            hd_data = (lhtx_tid_hold[7:6] == 2'b00) ? {40'bx,LA_lhtx_tdata[63:40]} : {56'bx,LA_lhtx_tdata[63:56]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = (lhtx_tid_hold[7:6] == 2'b00) ? 1'b0 : (!LA_lhtx_tkeep[6]);
            hd_we   = (lhtx_tid_hold[7:6] == 2'b00) ? 8'b0000_0111 : 8'b0000_0001;
            hd_vld  = 1'b1;
          end
          default: begin
            hd_keep = lhtx_tlast_hold ?  ((lhtx_tid_hold[7:6] == 2'b00) ? {lhtx_tkeep_hold[4:0],3'b0} : {lhtx_tkeep_hold[6:0],1'b0}) : 8'b1111_1111;
            hd_data = (lhtx_tid_hold[7:6] == 2'b00) ? {hello_data_hold[39:0],LA_lhtx_tdata[63:40]} : {hello_data_hold[55:0],LA_lhtx_tdata[63:56]};
            hd_user = 8'bxxxx_xxxx;
            hd_last =  (LA_lhtx_tlast & (((lhtx_tid_hold[7:6] == 2'b00) & (!LA_lhtx_tkeep[4])) || 
                       ((lhtx_tid_hold[7:6] != 2'b00) & (!LA_lhtx_tkeep[6])))) ? 1'b1 :  lhtx_tlast_hold ;
            hd_we   = hd_update ? 8'b1111_1111 : 8'b0000_0000;
            hd_vld  = hd_update;
       
          end
        endcase
      end
      default: begin
            hd_keep = 8'hFF;
            hd_data = 64'bx;
            hd_user = 8'bxxxx_xxxx;
            hd_last = 1'b0;
            hd_we   = 8'b0000_0000;
            hd_vld  = 1'b0;
      end
    endcase
  end
end // end if (DEVICEID_WIDTH == 8)
// When using 16-bit device IDs, data alignment is different
else begin: hello_decoder_16devid_gen // if (DEVICEID_WIDTH == 16)
  always @* begin
    case ({1'b0,lhtx_ftype})
      FTYPE_NREAD,FTYPE_NWRITE: begin
        case ({hd_first,hd_second})
          2'b10: begin
            hd_keep = 8'b1111_1111;
            hd_data = {hello_prio,TT,hello_ftype,hello_destid,hello_srcid,hello_ttype,
                       hello_rdwrsize,hello_tid,hello_addr[31:24]};
            hd_user = {3'b0,1'b0,1'b0,hello_vc,hello_crf,1'b0};
            hd_last = 1'b0;
            hd_we   = 8'b1111_1111;
            hd_vld  = 1'b1;
          end
          2'b01: begin
            hd_keep = lhtx_tlast_hold ? 8'b1110_0000 : 8'b1111_1111;
            hd_data = {hello_addr_hold[23:3],hello_wdptr_hold,hello_xamsbs_hold,LA_lhtx_tdata[63:24]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = lhtx_tlast_hold;
            hd_we   = 8'b1111_1111;
            hd_vld  = 1'b1;
          end
          default: begin
            hd_keep = lhtx_tlast_hold ? 8'b1110_0000 : 8'b1111_1111;
            hd_data = {hello_data_hold[23:0],LA_lhtx_tdata[63:24]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = lhtx_tlast_hold;
            hd_we   = hd_update ? 8'b1111_1111 : 8'b0000_0000;
            hd_vld  = hd_update;
          end
        endcase
      end
      FTYPE_SWRITE: begin
        case ({hd_first,hd_second})
          2'b10: begin
            hd_keep = 8'b1111_1111;
            hd_data = {hello_prio,TT,hello_ftype,hello_destid,hello_srcid,
                       hello_addr[31:8]};
            hd_user = {3'b0,1'b0,1'b0,hello_vc,hello_crf,1'b0};
            hd_last = 1'b0;
            hd_we   = 8'b1111_1111;
            hd_vld  = 1'b1;
          end
          2'b01: begin
            hd_keep = 8'b1111_1111;
            hd_data = {hello_addr_hold[7:3],1'b0,hello_xamsbs_hold,LA_lhtx_tdata[63:8]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = 1'b0;
            hd_we   = 8'b1111_1111;
            hd_vld  = 1'b1;
          end
          default: begin
            hd_keep = lhtx_tlast_hold ? 8'b1000_0000 : 8'b1111_1111;
            hd_data = {hello_data_hold[7:0],LA_lhtx_tdata[63:8]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = lhtx_tlast_hold;
            hd_we   = hd_update ? 8'b1111_1111 : 8'b0000_0000;
            hd_vld  = hd_update;
          end
        endcase
      end
      FTYPE_MAINT: begin
        case ({hd_first,hd_second})
          2'b10: begin
            hd_keep = 8'b1111_1111;
            hd_data = {hello_prio,TT,hello_ftype,hello_destid,hello_srcid,hello_ttype,
                       hello_sizestat,hello_tid,hello_addr[31:24]};
            hd_user = {3'b0,hello_maintresp,1'b0,hello_vc,hello_crf,1'b0};
            hd_last = 1'b0;
            hd_we   = 8'b1111_1111;
            hd_vld  = 1'b1;
          end
          2'b01: begin
            hd_keep = lhtx_tlast_hold ? 8'b1110_0000 : 8'b1111_1111;
            hd_data = {hello_addr_hold[23:3],hello_wdptr_hold,2'b0,LA_lhtx_tdata[63:24]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = lhtx_tlast_hold;
            hd_we   = 8'b1111_1111;
            hd_vld  = 1'b1;
          end
          default: begin
            hd_keep = lhtx_tlast_hold ? 8'b1110_0000 : 8'b1111_1111;
            hd_data = {hello_data_hold[23:0],LA_lhtx_tdata[63:24]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = lhtx_tlast_hold;
            hd_we   = hd_update ? 8'b1111_1111 : 8'b0000_0000;
            hd_vld  = hd_update;
          end
        endcase
      end
      FTYPE_MSG: begin
        case ({hd_first,hd_second})
          2'b10: begin
            hd_keep = 8'b1111_1111;
            hd_data = {hello_prio,TT,hello_ftype,hello_destid,hello_srcid,hello_msglen,
                       hello_ssize,hello_letter,hello_mbox,hello_msgsegxmbox,8'bx};
            hd_user = {3'b0,1'b0,1'b0,hello_vc,hello_crf,1'b0};
            hd_last = 1'b0;
            hd_we   = 8'b1111_1110;
            hd_vld  = 1'b0;
          end
          2'b01: begin
            hd_keep = 8'b1111_1111;
            hd_data = {56'bx,LA_lhtx_tdata[63:56]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = 1'b0;
            hd_we   = 8'b0000_0001;
            hd_vld  = 1'b1;
          end
          default: begin
            hd_keep = lhtx_tlast_hold ? 8'b1111_1110 : 8'b1111_1111;
            hd_data = {hello_data_hold[55:0],LA_lhtx_tdata[63:56]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = lhtx_tlast_hold;
            hd_we   = hd_update ? 8'b1111_1111 : 8'b0000_0000;
            hd_vld  = hd_update;
          end
        endcase
      end
      FTYPE_DB: begin
        case ({hd_first,hd_second})
          2'b10: begin
            hd_keep = 8'b1111_1111;
            hd_data = {hello_prio,TT,hello_ftype,hello_destid,hello_srcid,
                       8'b0,hello_tid,hello_addr[31:24]};
            hd_user = {3'b0,1'b0,1'b0,hello_vc,hello_crf,1'b0};
            hd_last = 1'b0;
            hd_we   = 8'b1111_1111;
            hd_vld  = 1'b1;
          end
          default: begin
            hd_keep = 8'b1000_0000;
            hd_data = {hello_addr_hold[23:16],56'bx};
            hd_user = 8'bxxxx_xxxx;
            hd_last = 1'b1;
            hd_we   = hd_update ? 8'b1000_0000 : 8'b0000_0000;
            hd_vld  = hd_update;
          end
        endcase
      end
      FTYPE_RESP: begin
        case ({hd_first,hd_second})
          2'b10: begin
            hd_keep = LA_lhtx_tlast ? 8'b1111_1110 : 8'b1111_1111;
            hd_data = {hello_prio,TT,hello_ftype,hello_destid,hello_srcid,hello_ttype,hello_stat,
                       hello_tid,8'bx};
            hd_user = {3'b0,1'b1,1'b0,hello_vc,hello_crf,1'b0};
            hd_last = LA_lhtx_tlast;
            hd_we   = 8'b1111_1110;
            hd_vld  = LA_lhtx_tlast;
          end
          2'b01: begin
            hd_keep = 8'b1111_1111;
            hd_data = {56'bx,LA_lhtx_tdata[63:56]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = 1'b0;
            hd_we   = 8'b0000_0001;
            hd_vld  = 1'b1;
          end
          default: begin
            hd_keep = lhtx_tlast_hold ? 8'b1111_1110 : 8'b1111_1111;
            hd_data = {hello_data_hold[55:0],LA_lhtx_tdata[63:56]};
            hd_user = 8'bxxxx_xxxx;
            hd_last = lhtx_tlast_hold;
            hd_we   = hd_update ? 8'b1111_1111 : 8'b0000_0000;
            hd_vld  = hd_update;
          end
        endcase
      end
      FTYPE_DS: begin
        case ({hd_first,hd_second})
          2'b10: begin
            hd_keep = 8'b1111_1111;
            hd_data = {hello_prio,TT,hello_ftype,hello_destid,hello_srcid,hello_size,
                       hello_tid,(hello_tid[7:6] == 2'b01 ? hello_addr[15:8] : hello_addr[31:24])};
            hd_user = {3'b0,1'b0,1'b0,hello_vc,hello_crf,1'b0};
            hd_last = 1'b0;
            hd_we   = (hello_tid[7:6] == 2'b00) ? 8'b1111_1110 : 8'b1111_1111;
            hd_vld  = (hello_tid[7:6] == 2'b00) ? 1'b0 : 1'b1;
          end
          2'b01: begin
            hd_keep =  (lhtx_tid_hold[7:6] == 2'b00) ? 8'b1111_1111 :
                       (LA_lhtx_tlast ? {1'b1,LA_lhtx_tkeep[7:1]} : 8'b1111_1111); 
            hd_data =  (lhtx_tid_hold[7:6] == 2'b00) ? 
                       {56'bx,LA_lhtx_tdata[63:56]} :
                       ({((lhtx_tid_hold[7:6] == 2'b01) ? hello_data_hold[7:0] : hello_data_hold[23:16]),
	               LA_lhtx_tdata[63:8]});
            hd_user = 8'bxxxx_xxxx;
            hd_last = (lhtx_tid_hold[7:6] == 2'b00) ? 1'b0 : (!LA_lhtx_tkeep[0]);
            hd_we   = hd_update ? ((lhtx_tid_hold[7:6] == 2'b00) ? 8'b0000_0001 : 8'b1111_1111) : 8'b0000_0000;
            hd_vld  = hd_update;
          end
          default: begin
       
            hd_keep = lhtx_tlast_hold ?  ((lhtx_tid_hold[7:6] == 2'b00) ? {lhtx_tkeep_hold[6:0],1'b0} : {lhtx_tkeep_hold[0],7'b0}) :
	              ((lhtx_tid_hold[7:6] == 2'b00) ? {lhtx_tkeep_hold[6:0],LA_lhtx_tkeep[7]} : {lhtx_tkeep_hold[0],LA_lhtx_tkeep[7:1]});

            hd_data = (lhtx_tid_hold[7:6] == 2'b00) ? {hello_data_hold[55:0],LA_lhtx_tdata[63:56]} : {hello_data_hold[7:0],LA_lhtx_tdata[63:8]};
            hd_user = 8'bxxxx_xxxx;
            hd_last =  (LA_lhtx_tlast & hd_update & (((lhtx_tid_hold[7:6] == 2'b00) & (!LA_lhtx_tkeep[6] )) || 
                       ((lhtx_tid_hold[7:6] != 2'b00) & (!LA_lhtx_tkeep[0])))) ? 1'b1 :  lhtx_tlast_hold;
            hd_we   = hd_update ? 8'b1111_1111 : 8'b0000_0000;
            hd_vld  = hd_update;
          
          end
        endcase
      end
      default: begin
            hd_keep = 8'hFF;
            hd_data = 64'bx;
            hd_user = 8'bxxxx_xxxx;
            hd_last = 1'b0;
            hd_we   = 8'b0000_0000;
            hd_vld  = 1'b0;
      end
    endcase
  end
end endgenerate // end if (DEVICEID_WIDTH == 16)

  // Decode FTYPE and TTYPE so that the RESPONSE bit of TUSER can be set appropriately
  // These signals are only valid on lhtx_sof
  assign srio_ftype = LA_lhtx_tdata[3:0];
  assign srio_ttype = (DEVICEID_WIDTH == 8) ? LA_lhtx_tdata[31:28] : LA_lhtx_tdata[47:44];
  assign srio_resp  = ((srio_ftype ==  FTYPE_RESP[3:0]) ||
                       (srio_ftype == FTYPE_MAINT[3:0]) && (srio_ttype[3:1] == 3'b001));

  // Re-swizzle decoded packet before sending to buffer
  assign bn_data   = {hd_data[7:0],   hd_data[15:8],  hd_data[23:16], hd_data[31:24],
                      hd_data[39:32], hd_data[47:40], hd_data[55:48], hd_data[63:56]};
  assign bn_keep   = {hd_keep[0],     hd_keep[1],     hd_keep[2],     hd_keep[3],
                      hd_keep[4],     hd_keep[5],     hd_keep[6],     hd_keep[7]};
  assign bn_we     = {hd_we[0],       hd_we[1],       hd_we[2],       hd_we[3],
                      hd_we[4],       hd_we[5],       hd_we[6],       hd_we[7]};

  // Mux between the decoded packet and the input data based on whether the packet uses HELLO format
  assign buft_keep = !hello_decode ? LA_lhtx_tkeep : bn_keep;
  assign buft_data =  hello_decode ? bn_data :  LA_lhtx_tdata;
  assign buft_we   =  hello_decode ? bn_we   :  8'hFF;
  assign buft_user =  hello_decode ? hd_user : {LA_lhtx_tuser[7:5], srio_resp, LA_lhtx_tuser[3:0]};
  assign buft_last =  hello_decode ? hd_last :  LA_lhtx_tlast;
  assign buft_vld  =  hello_decode ? hd_vld  :  lhtx_active;

  //*ASSERTION*
  //(ap_not_lhtx_second_and_lhtx_sof): lhtx_second should not be asserted on lhtx_sof

  // }}} Create sRIO Native packet

  //Register the keep, data, and user bits so they're available if the buffer stalls
  always @(posedge log_clk) begin
    // No reset needed because only sampled on valid
    if (buffer_stall && !buffer_stall_q) begin
      if (lhtx_sof) begin
        holdreg_tuser <= #TCQ buft_user;
      end
      holdreg_tkeep   <= #TCQ buft_keep;
      // Only write the data bytes that are enabled (this saves registers)
      if (buft_we[7])
        holdreg_tdata[63:56] <= #TCQ buft_data[63:56];
      if (buft_we[6])
        holdreg_tdata[55:48] <= #TCQ buft_data[55:48];
      if (buft_we[5])
        holdreg_tdata[47:40] <= #TCQ buft_data[47:40];
      if (buft_we[4])
        holdreg_tdata[39:32] <= #TCQ buft_data[39:32];
      if (buft_we[3])
        holdreg_tdata[31:24] <= #TCQ buft_data[31:24];
      if (buft_we[2])
        holdreg_tdata[23:16] <= #TCQ buft_data[23:16];
      if (buft_we[1])
        holdreg_tdata[15:8]  <= #TCQ buft_data[15:8];
      if (buft_we[0])
        holdreg_tdata[7:0]   <= #TCQ buft_data[7:0];
    end
  end

  // {{{ Output Generation
  // + {{{ Buffer Interface +

  // Register the keep, data, and user bits for the output
  // After a buffer stall, grab data from holdreg, otherwise directly from mux
  always @(posedge log_clk) begin
    // No reset needed because only sampled on valid
    if (!buffer_stall) begin
      if (buffer_stall_fell && buffer_stall_active) begin
        LD_buft_tkeep <= #TCQ holdreg_tkeep;
        LD_buft_tdata <= #TCQ holdreg_tdata;
        if (buffer_stall_sof) begin
          LD_buft_tuser <= #TCQ holdreg_tuser;
        end
      end else begin
        if (lhtx_sof) begin
          LD_buft_tuser <= #TCQ buft_user;
        end
        LD_buft_tkeep <= #TCQ buft_keep;
        //Only write the data bytes that are enabled (this saves registers)
        if (buft_we[7])
          LD_buft_tdata[63:56] <= #TCQ buft_data[63:56];
        if (buft_we[6])
          LD_buft_tdata[55:48] <= #TCQ buft_data[55:48];
        if (buft_we[5])
          LD_buft_tdata[47:40] <= #TCQ buft_data[47:40];
        if (buft_we[4])
          LD_buft_tdata[39:32] <= #TCQ buft_data[39:32];
        if (buft_we[3])
          LD_buft_tdata[31:24] <= #TCQ buft_data[31:24];
        if (buft_we[2])
          LD_buft_tdata[23:16] <= #TCQ buft_data[23:16];
        if (buft_we[1])
          LD_buft_tdata[15:8]  <= #TCQ buft_data[15:8];
        if (buft_we[0])
          LD_buft_tdata[7:0]   <= #TCQ buft_data[7:0];
      end
    end
  end

  // Create TLAST - during stall - hold value, after a stall - look at holdreg, else use mux value
  assign ld_buft_tlast_d  = (buffer_stall_fell) ? buffer_stall_last :
                            !buffer_stall ? buft_last : LD_buft_tlast;
  // Create TVALID - during stall - hold value, after a stall - look at value before stall,
  //                 else use mux value plus indicate valid if a beat is supposed to be inserted
  assign ld_buft_tvalid_d = buffer_stall        ? LD_buft_tvalid :
                            buffer_stall_fell   ? buffer_stall_valid :
                            buffer_stall_fell_q && hd_insert_beat || ((lhtx_active || hd_insert_beat) && buft_vld);

  // Register TLAST and TVALID
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LD_buft_tvalid <= #TCQ 1'b0;
      LD_buft_tlast  <= #TCQ 1'b0;
    end else begin
      LD_buft_tvalid <= #TCQ ld_buft_tvalid_d;
      LD_buft_tlast  <= #TCQ ld_buft_tlast_d;
    end
  end


  // Internal Coverage and Assertions
  //*COVERAGE*
  //(cp_partial_write_of_buft_data): Only some of the data bytes are written

  // Buffer Interface Coverage and Assertions
  //*COVERAGE*
  //(cp_tx_rb2b_two_single_cycle_pkts): cover that back to back single cycle packets exit the buffer
  //(cp_buft_buffer_stalls_mid_packet): The buffer stalls mid-packet
  //(cp_buft_buffer_stalls_btw_packets): The buffer stalls between packets
  //(cp_buft_buffer_stalls_first_beat): The buffer stalls after the first beat

  //*ASSERTION*
  //(ap_buft_valid_high_until_active): Once asserted, LD_buft_tvalid stays high until BT_buft_tready is asserted

  // + }}} end Buffer Interface +

  // + {{{ Arbiter Interface +

  // Create the TREADY signal for the lhtx interface
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LD_lhtx_tready <= #TCQ 1'b0;
    end else begin
      LD_lhtx_tready <= #TCQ !(buffer_stall ||                       // Backpressure if buffer stalls
                               need_extra_beat ||                    // or if an extra beat is required b/c of HELLO
                               buffer_stall_fell && hd_insert_beat); // or if there's an extra beat req during stall
    end
  end

  // Arbiter Interface Coverage and Assertions
  //*COVERAGE*
  //(cp_lhtx_b2b_single_cycle): There are back-to-back single-cycle packets on the lhtx interface
  //(cp_lhtx_arbiter_stalls_mid_packet): The arbiter stalls mid-packet
  //(cp_lhtx_arbiter_stalls_btw_packets): The arbiter stalls between packets
  //(cp_lhtx_arbiter_stalls_first_beat): The arbiter stalls after the first beat
  //(cp_lhtx_hd_stalls_mid_packet): The hello_decoder stalls mid-packet
  //(cp_lhtx_hd_stalls_btw_packets): The hello_decoder stalls between packets
  //(cp_lhtx_hd_stalls_first_beat): The hello_decoder stalls after the first beat

  //*ASSERTION*
  //(ap_lhtx_valid_high_until_active): Once asserted, LA_lhtx_tvalid stays high until LD_lhtx_tready is asserted
  //(ap_lhtx_hello_tkeep_all_ones): LA_lhtx_tkeep is 8'hFF on valid cycles of HELLO packets

  // + }}} end Arbiter Interface +
  // }}} Output Generation


endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/log/log_cfg/srio_gen2_v4_1_16_log_cfg_reg.v#2 $
//----------------------------------------------------------------------
//
// LOG_CFG_REG
// Description:
// This module contains the configuration registers for the LOG layer.
//
// For writes, it takes a write enable, address, data and strobe (byte
// enables) from the cfg_axi module and handles writes to writable
// registers. For reads, it takes an address and read enable, and
// returns the read data from the corresponding CSR. It also has a LOG
// core interface for transfer of control and status information.
//
// To view the CSR in simulation, pull the csr_log_xxx wire.
//
// Hierarchy:
// LOG_TOP
//    |______LOG_CFG_TOP
//              |______CFG_AXI (in hdl/common/)
//              |______LOG_CFG_REG <-- this module
// ---------------------------------------------------------------------
`timescale 1ps/1ps

module srio_gen2_v4_1_16_log_cfg_reg
  #(
    parameter TCQ             = 100,
    parameter HW_ARCH         = 2,        // Device {V5LXT(0), V5FXT(1), V6LXT(2), V6CXT(3), S6LXT(4)}
    parameter DEVICEID_WIDTH  = 8,        // Source/Destination ID width {8,16}
    parameter DEVICEID        = 16'h00FF, // Reset value for Device ID {16'h0000-16'hFFFF}
    parameter INIT_NREAD      = 1,        // Core may initiate NREAD transactions {0,1}
    parameter INIT_NWRITE     = 1,        // Core may initiate NWRITE transactions {0,1}
    parameter INIT_SWRITE     = 1,        // Core may initiate SWRITE transactions {0,1}
    parameter INIT_NWRITE_R   = 1,        // Core may initiate NWRITE_R transactions {0,1}
    parameter INIT_DB         = 1,        // Core may initiate Doorbell transactions {0,1}
    parameter INIT_DS         = 1,        // Core may initiate Data-Streaming transactions {0,1}
    parameter INIT_ATOMIC     = 1,        // Core may initiate ATOMIC transactions {0,1}
    parameter MSG_INIT_SINGLE = 1,        // Core may initiate single-segment message transactions {0,1}
    parameter MSG_INIT_MULTI  = 1,        // Core may initiate multiple-segment message transactions {0,1}
    parameter TARGET_NREAD    = 1,        // Core may sink NREAD transactions {0,1}
    parameter TARGET_NWRITE   = 1,        // Core may sink NWRITE transactions {0,1}
    parameter TARGET_SWRITE   = 1,        // Core may sink SWRITE transactions {0,1}
    parameter TARGET_NWRITE_R = 1,        // Core may sink NWRITE_R transactions {0,1}
    parameter TARGET_DB       = 1,        // Core may sink Doorbell transactions {0,1}
    parameter TARGET_DS       = 1,        // Core may sink Data-Streaming transactions {0,1}
    parameter TARGET_ATOMIC   = 1,        // Core may sink ATOMIC transactions {0,1}
    parameter MSG_SINK_SINGLE = 1,        // Core may sink single-segment message transactions {0,1}
    parameter MSG_SINK_MULTI  = 1,        // Core may sink multiple-segment message transactions {0,1}
    parameter CRF_SUPPORT     = 1,        // If set, the core supports use of the CRF flag {0,1}
    parameter DEVID_CAR       = 32'h00000000, // Reset value for Device Identity CAR {32�h00000000�?32�hFFFFFFFF}
    parameter DEVINFO_CAR     = 32'h00000000, // Reset value for Device Info CAR {32�h00000000�?32�hFFFFFFFF}
    parameter DEV_CAR_OVRD    = 0,            // If 1, DEV*CAR param values used {0,1}
    parameter LCSBA_SUPPORT   = 1,        // If set, the LCSBA is used to reroute transactions to the maint port {0,1}
    parameter LCSBA           = 10'h3FF,  // Reset value for LCSBA register {10'h0-10'h3FF}
    parameter ASSY_ID         = 16'h0000, // Assembly ID from GUI {16'h0000-16'hFFFF}
    parameter ASSY_VENDOR     = 16'h0000, // Assembly Vendor ID from GUI {16'h0000-16'hFFFF}
    parameter ASSY_REV        = 16'h0000, // Assembly Revision from GUI {16'h0000-16'hFFFF}
    parameter PE_BRIDGE       = 0,        // Processing Element contains Bridge functionality {0,1}
    parameter PE_MEMORY       = 1,        // Processing Element contains Memory functionality {0,1}
    parameter PE_PROC         = 0,        // Processing Element contains Processor functionality {0,1}
    parameter PE_SWITCH       = 0,        // Processing Element contains Switch functionality {0,1}
    parameter PHY_EF_PTR      = 16'h0100  // Location of PHY ext features {0x0100+}
  )(
    // {{{ Port Declarations ---------------
    // System Signals
    input             log_clk,                  // LOG interface clock
    input             log_rst,                  // Reset for LOG clock Domain
    input             CCA_sync_cfg_rst,         // cfg_rst sync'ed to log_clk

    // User Interface
    // Current Device ID - Used as SourceID for transmitted packets
    output reg [15:0] LCR_deviceid = (DEVICEID_WIDTH == 8) ? {8'b0, DEVICEID[7:0]} : DEVICEID,

    // LOG Arb Interface
    output reg [9:0]  LCR_lcsba = LCSBA,        // Local Configuration Base Address register mask value

    // Generic Configuration Interface (cfg_axi sub-module)
    input      [23:0] CCA_cfg_waddr,            // Write Address
    input      [31:0] CCA_cfg_wdata,            // Write Data
    input      [3:0]  CCA_cfg_wstrb,            // Write Data Byte Enables
    input             CCA_sync_we,              // Synchronized write enable
    input      [23:0] CCA_cfg_raddr,            // Read Address
    input             CCA_sync_re,              // Synchronized Read Enable
    output reg [31:0] LCR_core_rdata            // Read Data
    // }}} End Port Declarations -----------
  );

// added below macro to fix the CR# 735137
// synthesis translate_off 
// {{{ Catch Bad Parameters
  //Catch any invalid parameter conditions
  initial begin
    //If the Device Identity Register does not have a value defined for the selected device, finish
    if ((HW_ARCH < 0) || (HW_ARCH > 14)) begin
      $display("ERROR: Invalid device selected for the LOG based on HW_ARCH=%0d.",
                HW_ARCH);
      $finish;
    end
  end
  // }}}
// synthesis translate_on 

  // {{{ Localparams -----------------------
  localparam        MAJOR_REV   =  4'h4;                    // Core Major Revision
  localparam        MINOR_REV   =  4'h0;                    // Core Minor Revision
  localparam        PATCH_REV   =  4'h0;                    // Core Patch Revision
  localparam        SPEC_REV    =  4'h2;                    // RapidIO Specification Revision (4'h2 indicates rev2.1)
  localparam        VENDORID    =  16'h000E;                // RIOTA-assigned Vendor ID
  localparam [3:0]  FAMILY      =  (HW_ARCH == 0) ? 4'h3 :  // Virtex (V5LXT)
                                   (HW_ARCH == 1) ? 4'h3 :  // Virtex (V5FXT)
                                   (HW_ARCH == 2) ? 4'h3 :  // Virtex (V6LXT)
                                   (HW_ARCH == 3) ? 4'h3 :  // Virtex (V6CXT)
                                   (HW_ARCH == 4) ? 4'h0 :  // Spartan (S6LXT)
                                   (HW_ARCH == 5) ? 4'h1 :  // Artix (A7T)
                                   (HW_ARCH == 6) ? 4'h2 :  // Kintex (K7T)
                                   (HW_ARCH == 7) ? 4'h3 :  // Virtex (V7T)
                                   (HW_ARCH == 8) ? 4'h3 :  // Virtex (V7XT)
                                   (HW_ARCH == 9) ? 4'h4 :  // Zynq
                                   (HW_ARCH == 10) ? 4'h2 :  // Ultrascale// this 2 is for KU devices
                                   (HW_ARCH == 11) ? 4'h3 :  // Ultrascale// this 3 is for VU devices
                                   (HW_ARCH == 12) ? 4'h4 :  // Ultrascale// this 4 is for ZUP devices
                                   (HW_ARCH == 13) ? 4'h5 :  // Ultrascale// this 5 is for KUP devices
                                   (HW_ARCH == 14) ? 4'h6 :  // Ultrascale// TBD alagarr
                                                    4'hF ;  // Default (undefined)

  localparam [3:0]  GENERATION  =  (HW_ARCH == 0) ? 4'h5 :  // 5 (V5LXT)
                                   (HW_ARCH == 1) ? 4'h5 :  // 5 (V5FXT)
                                   (HW_ARCH == 2) ? 4'h6 :  // 6 (V6LXT)
                                   (HW_ARCH == 3) ? 4'h6 :  // 6 (V6CXT)
                                   (HW_ARCH == 4) ? 4'h6 :  // 6 (S6LXT)
                                   (HW_ARCH == 5) ? 4'h7 :  // 7 (A7T)
                                   (HW_ARCH == 6) ? 4'h7 :  // 7 (K7T)
                                   (HW_ARCH == 7) ? 4'h7 :  // 7 (V7T)
                                   (HW_ARCH == 8) ? 4'h7 :  // 7 (V7XT)
                                   (HW_ARCH == 9) ? 4'h8 :  // 8 (Zynq)
                                   (HW_ARCH == 10) ? 4'h8 :  // 8 (Ultrascale)// both for ku and vu the no. 8 is same
                                   (HW_ARCH == 11) ? 4'h8 :  // 8 (Ultrascale)// both for ku and vu the no. 8 is same
                                   (HW_ARCH == 12) ? 4'h8 :  // 8 (Ultrascale)// both for ku and vu the no. 8 is same
                                   (HW_ARCH == 13) ? 4'h8 :  // 8 (Ultrascale)// both for ku and vu the no. 8 is same
                                   (HW_ARCH == 14) ? 4'h8 :  // 8 (Ultrascale)// both for ku and vu the no. 8 is same
                                                    4'hF ;  // Default (undefined)

  localparam [3:0]  LAST_VAL  =  (HW_ARCH == 10) ? 4'h5 : // this is added to make the KU or VU to appear as 
                                 (HW_ARCH == 11) ? 4'h5 : // 285 or 385
                                 (HW_ARCH == 12) ? 4'h5 : // 485
                                 (HW_ARCH == 13) ? 4'h5 : // 585
                                 (HW_ARCH == 14) ? 4'h5 : // 685
				                   4'h0;  // this is for non KU/VU devices

  localparam        INIT_MSG    =  MSG_INIT_SINGLE ||       // Core can initiate message transactions
                                   MSG_INIT_MULTI;

  localparam        TARGET_MSG  =  MSG_SINK_SINGLE ||       // Core can sink message transactions
                                   MSG_SINK_MULTI;


  // Parameters for CAR/CSR offsets
  // Capability Registers:
  localparam [15:0] LOG_000   =  16'h0000;  // Device Identity CAR
  localparam [15:0] LOG_004   =  16'h0004;  // Device Information CAR
  localparam [15:0] LOG_008   =  16'h0008;  // Assembly Identity CAR
  localparam [15:0] LOG_00C   =  16'h000C;  // Assembly Information CAR
  localparam [15:0] LOG_010   =  16'h0010;  // Processing Element Features CAR
  localparam [15:0] LOG_014   =  16'h0014;  // Switch Port Information CAR
  localparam [15:0] LOG_018   =  16'h0018;  // Source Operations CAR
  localparam [15:0] LOG_01C   =  16'h001C;  // Destination Operations CAR
  // Command and Status Registers:
  localparam [15:0] LOG_04C   =  16'h004C;  // Processing Element Logical Layer CSR
  localparam [15:0] LOG_058   =  16'h0058;  // Local Configuration Space High Base Address CSR
  localparam [15:0] LOG_05C   =  16'h005C;  // Local Configuration Space Base Address CSR
  localparam [15:0] LOG_060   =  16'h0060;  // Base Device ID CSR
  localparam [15:0] LOG_068   =  16'h0068;  // Host Base Device ID Lock CSR
  localparam [15:0] LOG_06C   =  16'h006C;  // Component Tag CSR
  // }}} End Localparams -------------------

  // {{{ Wire Declarations -----------------
                                                // placeholder for registered version of log_rst (currently not used)
  reg   [7:0]   base_deviceid = DEVICEID[7:0];  // Base_deviceID field for Base Device ID CSR
  reg   [15:0]  large_base_deviceid = DEVICEID; // Large_base_deviceID field for Base Device ID CSR
  reg   [15:0]  host_base_deviceid;             // Host_base_deviceID field for Host Base Device ID Lock CSR
  reg   [9:0]   writable_lcsba = LCSBA;         // Local Configuration Space Base Address from writable register
  reg   [31:0]  component_tag;                  // Component Tag field for Component Tag CSR
                // CSR is being written
  wire          log_05c_write, log_060_write, log_068_write, log_06c_write;
                // Assembled CSRs for easy simulation viewing
  wire  [31:0]  csr_log_000, csr_log_004, csr_log_008, csr_log_00c, csr_log_010,
                csr_log_014, csr_log_018, csr_log_01c, csr_log_04c, csr_log_058,
                csr_log_05c, csr_log_060, csr_log_068, csr_log_06c;

  // }}} End Wire Declarations -------------


  // {{{ Writable Register Bank ------------
  // A shadow register is kept for writable registers so that read and write
  // functionality can be fully separated.

  // Create signal to indicate that a given register is targeted for a write operation.
  // Only need to do this for registers with writable fields.
  assign log_05c_write = CCA_sync_we && (CCA_cfg_waddr[15:0] == LOG_05C);
  assign log_060_write = CCA_sync_we && (CCA_cfg_waddr[15:0] == LOG_060);
  assign log_068_write = CCA_sync_we && (CCA_cfg_waddr[15:0] == LOG_068);
  assign log_06c_write = CCA_sync_we && (CCA_cfg_waddr[15:0] == LOG_06C);


  // --------------- Command and Status Registers ------------------------
  // ----- Local Configuration Space Base Address CSR writable registers ----- //
  always @(posedge log_clk) begin
    if (CCA_sync_cfg_rst) begin
      writable_lcsba              <= #TCQ LCSBA[9:0];
    end else if (log_05c_write) begin
      if (CCA_cfg_wstrb[3])
        writable_lcsba[9:3]       <= #TCQ CCA_cfg_wdata[30:24];
      if (CCA_cfg_wstrb[2])
        writable_lcsba[2:0]       <= #TCQ CCA_cfg_wdata[23:21];
    end
  end

  // Create LCSBA output
  always @* begin
    LCR_lcsba = (LCSBA_SUPPORT == 1) ? writable_lcsba : LCSBA;
  end

  // ----- Base Device ID CSR writable registers ----- //
  always @(posedge log_clk) begin
    if (CCA_sync_cfg_rst) begin
      base_deviceid               <= #TCQ DEVICEID[7:0];
      large_base_deviceid         <= #TCQ DEVICEID[15:0];
    end else if (log_060_write) begin
      if (CCA_cfg_wstrb[2])
        base_deviceid[7:0]        <= #TCQ CCA_cfg_wdata[23:16];
      if (CCA_cfg_wstrb[1])
        large_base_deviceid[15:8] <= #TCQ CCA_cfg_wdata[15:8];
      if (CCA_cfg_wstrb[0])
        large_base_deviceid[7:0]  <= #TCQ CCA_cfg_wdata[7:0];
    end
  end

  // Create Device ID output
  always @* begin
    LCR_deviceid = (DEVICEID_WIDTH == 8) ? {8'b0, base_deviceid} : large_base_deviceid;
  end

  // ----- Host Base Device ID Lock CSR writable registers ----- //
  // The Host_base_deviceID field is write-once/resetable with a lock function.
  // Once the Host_base_deviceID field is written, subsequent writes are
  // ignored unless the value written matches the value stored in the field, in
  // which case the register is re-initialized to 16'hFFFF
  always @(posedge log_clk) begin
    if (CCA_sync_cfg_rst) begin
      host_base_deviceid          <= #TCQ 16'hFFFF;
    end else if (log_068_write) begin
      if (CCA_cfg_wstrb[1:0] == 2'b11) begin  // Only process write if both bytes are enabled
        if (host_base_deviceid == 16'hffff) begin
          // If Host_base_deviceID is 16'hFFFF, capture new value
          host_base_deviceid      <= #TCQ CCA_cfg_wdata[15:0];
        end else if (host_base_deviceid == CCA_cfg_wdata[15:0]) begin
          // If Host_base_deviceID is equal to the write value, reset to 16'hFFFF
          host_base_deviceid        <= #TCQ 16'hffff;
        end
      end
    end
  end

  //*COVERGROUP*
  //(cg_host_base_deviceid_enum): Enumerate host_base_deviceid field in Host Base Device ID Lock CSR

  //*ASSERTION*
  //(ap_host_base_deviceid_unlocks): The Host Base Device ID Lock CSR unlocks when written with stored value

  //*COVERPOINT*
  //(cp_unlock_host_base_deviceid): The Host Base Device ID Lock CSR is written with
  // the value stored in the CSR while the CSR is locked

  //*ASSERTION*
  //(ap_host_base_deviceid_updates_when_unlocked): Host_base_deviceID takes on the written value when unlocked

  //*COVERPOINT*
  //(cp_write_host_base_deviceid_with_ffff_value_when_not_locked): A write of 16'hFFF is received while
  // the Host Base Device ID Lock CSR is not locked

  //*COVERPOINT*
  //(cp_write_host_base_deviceid_with_other_value_when_not_locked): A write of !16'hFFFF is received while
  // the Host Base Device ID Lock CSR is not locked

  //*ASSERTION*
  //(ap_host_base_deviceid_ignores_partial_write): Host_base_deviceID does not change unless both bytes are written

  //*COVERGROUP*
  //(cg_host_base_deviceid_strb): Enumerate strobe for write to Host Base Device ID Lock CSR (host_base_deviceid field)

  //*ASSERTION*
  //(ap_host_base_deviceid_ignores_write_when_locked): Host_base_deviceID does not change when locked

  //*COVERPOINT*
  //(cp_write_log_068_when_locked): A write is received while the Host Base Device ID Lock CSR is locked

  //*COVERPOINT*
  //(cp_write_log_068_with_nonlock_value_when_locked): The Host Base Device ID Lock CSR is written with
  // a value not stored in the CSR while the CSR is locked

  // ----- Component Tag CSR writable registers ----- //
  always @(posedge log_clk) begin
    if (CCA_sync_cfg_rst) begin
      component_tag             <= #TCQ 32'b0;
    end else if (log_06c_write) begin
      if (CCA_cfg_wstrb[3])
        component_tag[31:24]    <= #TCQ CCA_cfg_wdata[31:24];
      if (CCA_cfg_wstrb[2])
        component_tag[23:16]    <= #TCQ CCA_cfg_wdata[23:16];
      if (CCA_cfg_wstrb[1])
        component_tag[15:8]     <= #TCQ CCA_cfg_wdata[15:8];
      if (CCA_cfg_wstrb[0])
        component_tag[7:0]      <= #TCQ CCA_cfg_wdata[7:0];
    end
  end
  // }}} End Writable Register Bank ---------

  // {{{ Read Data Assembly ----------------
  // Form read data based on address
  // Bit ordering mirrors RapidIO Spec (e.g. spec bit 0 -> log_cfg bit 31)

  // Create wires for each CAR/CSR for easy simulation viewing.
  // -------------------- Capability Registers ------------------------------------
                                                    // core  (spec)   Description
                                                    // ----------------------------
  // Device Identity CAR
  assign csr_log_000 = DEV_CAR_OVRD ? DEVID_CAR :   // 31:0   (0:31)  User override value
                       {4'b0,                       // 31:28  (0:3)   DeviceIdentity - reserved
                        FAMILY,                     // 27:24  (4:7)   DeviceIdentity - Family
                        GENERATION,                 // 23:20  (8:11)  DeviceIdentity - Generation
                        //4'b0,                       // 19:16  (12:15) DeviceIdentity - reserved
			LAST_VAL,            
                        VENDORID};                  // 15:0   (16:31) DeviceVendorIdentity

  // Device Information CAR
  assign csr_log_004 = DEV_CAR_OVRD ? DEVINFO_CAR : // 31:0   (0:31)  User override value
                       {12'b0,                      // 31:20  (0:11)  DeviceRev - reserved
                        SPEC_REV,                   // 19:16  (12:15) DeviceRev - Spec Revision (4'h2 indicates rev2.1)
                        4'b0,                       // 15:12  (16:19) DeviceRev - reserved
                        MAJOR_REV,                  // 11:8   (20:23) DeviceRev - Core Major Revision
                        MINOR_REV,                  // 7:4    (24:27) DeviceRev - Core Minor Revision
                        PATCH_REV};                 // 3:0    (28:31) DeviceRev - Core Patch Revision

  // Assembly Identity CAR
  assign csr_log_008 = {ASSY_ID[15:0],              // 31:16  (0:15)  AssyIdentity
                        ASSY_VENDOR[15:0]};         // 15:0   (16:31) AssyVendorIdentity

  // Assembly Information CAR
  assign csr_log_00c = {ASSY_REV[15:0],             // 31:16  (0:15)  AssyRev
                        PHY_EF_PTR[15:0]};          // 15:0   (16:31) ExtendedFeaturesPtr

  // Processing Element Features CAR
  assign csr_log_010 = {(PE_BRIDGE == 1),           // 31     (0)     Bridge
                        (PE_MEMORY == 1),           // 30     (1)     Memory
                        (PE_PROC == 1),             // 29     (2)     Processor
                        (PE_SWITCH == 1),           // 28     (3)     Switch
                        1'b0,                       // 27     (4)     Multiport
                        21'b0,                      // 26:4   (5:25)  Reserved, Implementation-defined
                        (CRF_SUPPORT == 1),         // 5      (26)    CRF support
                        (DEVICEID_WIDTH == 16),     // 4      (27)    Device ID Width 
                        1'b1,                       // 3      (28)    Extended features
                        3'b001};                    // 2:0    (29:31) Extended addressing support

  //FIXSWITCH Switch Port Information CAR - Placeholder, not valid if not a switch.
  assign csr_log_014 = {16'b0,                      // 31:16  (0:15)  Reserved
                        8'h00,                      // 15:8   (16:23) PortTotal
                        8'h00};                     // 7:0    (24:31) PortNumber

  // Source Operations CAR
  assign csr_log_018 = {13'b0,                      // 31:19  (0:12)  Reserved, Implementation Defined
                        (INIT_DS == 1),             // 18     (13)    Data-Streaming
			2'b0,                       // 17:16  (14:15) Implementation Defined
                        (INIT_NREAD == 1),          // 15     (16)    Read
                        (INIT_NWRITE == 1),         // 14     (17)    Write
                        (INIT_SWRITE == 1),         // 13     (18)    Streaming-write
                        (INIT_NWRITE_R == 1),       // 12     (19)    Write-with-response
                        (INIT_MSG == 1),            // 11     (20)    Data message
                        (INIT_DB == 1),             // 10     (21)    Doorbell
                        (INIT_ATOMIC == 1),         // 9      (22)    Atomic (compare-and-swap)
                        (INIT_ATOMIC == 1),         // 8      (23)    Atomic (test-and-swap)
                        (INIT_ATOMIC == 1),         // 7      (24)    Atomic (increment)
                        (INIT_ATOMIC == 1),         // 6      (25)    Atomic (decrement)
                        (INIT_ATOMIC == 1),         // 5      (26)    Atomic (set)
                        (INIT_ATOMIC == 1),         // 4      (27)    Atomic (clear)
                        (INIT_ATOMIC == 1),         // 3      (28)    Atomic (swap)
                        1'b0,                       // 2      (29)    Port-write
                        2'b0};                      // 1:0    (30:31) Implementation Defined

  // Destination Operations CAR
  assign csr_log_01c = {13'b0,                      // 31:19  (0:12)  Reserved, Implementation Defined
                        (TARGET_DS == 1),           // 18     (13)    Data-Streaming
			2'b0,                       // 17:16  (14:15) Implementation Defined
                        (TARGET_NREAD == 1),        // 15     (16)    Read
                        (TARGET_NWRITE == 1),       // 14     (17)    Write
                        (TARGET_SWRITE == 1),       // 13     (18)    Streaming-write
                        (TARGET_NWRITE_R == 1),     // 12     (19)    Write-with-response
                        (TARGET_MSG == 1),          // 11     (20)    Data message
                        (TARGET_DB == 1),           // 10     (21)    Doorbell
                        (TARGET_ATOMIC == 1),       // 9      (22)    Atomic (compare-and-swap)
                        (TARGET_ATOMIC == 1),       // 8      (23)    Atomic (test-and-swap)
                        (TARGET_ATOMIC == 1),       // 7      (24)    Atomic (increment)
                        (TARGET_ATOMIC == 1),       // 6      (25)    Atomic (decrement)
                        (TARGET_ATOMIC == 1),       // 5      (26)    Atomic (set)
                        (TARGET_ATOMIC == 1),       // 4      (27)    Atomic (clear)
                        (TARGET_ATOMIC == 1),       // 3      (28)    Atomic (swap)
                        1'b0,                       // 2      (29)    Port-write
                        2'b0};                      // 1:0    (30:31) Implementation Defined

  // -------------------- Command and Status Registers ----------------------------
                                                    // core  (spec)   Description
                                                    // ----------------------------
  // Processing Element Logical Layer CSR
  assign csr_log_04c = {29'b0,                      // 31:3   (0:28)  Reserved
                        3'b001};                    // 2:0    (29:31) Extended addressing control

  // Local Configuration Space Base Address 0 CSR
  assign csr_log_058 = {32'b0};                     // 31:0   (0:31)  Reserved for 34-bit local physical address

  // Local Configuration Space Base Address 1 CSR
  assign csr_log_05c = {1'b0,                       // 31     (0)     Reserved for 34-bit local physical address
                        LCR_lcsba, 21'b0};          // 30:0   (1:31)  LCSBA

  // Base Device ID CSR
  assign csr_log_060 = {8'b0,                       // 31:24  (0:7)   Reserved
                        base_deviceid,              // 23:16  (8:15)  Large_base_deviceID
                        large_base_deviceid};       // 15:0   (16:31) Large_base_deviceID

  // Host Base Device ID Lock CSR
  assign csr_log_068 = {16'b0,                      // 31:16  (0:15)  Reserved
                        host_base_deviceid};        // 15:0   (16:31) Host_base_deviceID

  // Component Tag CSR
  assign csr_log_06c = component_tag;               // 31:0   (0:31)  component_tag

  //*COVERAGE*
  //(cp_log_000_rd_b4_wr): Cover that each byte of log_000 was read before it was written
  //(cp_log_000_rd_aftr_wr): Cover that each byte of log_000 was read after it was written
  //(cp_log_000_3_rst_val_chk): Cover that HW_ARCH is non-default and log_000 byte 3 was rd_b4_wr
  //(cp_log_000_2_rst_val_chk): Cover that HW_ARCH is non-default and log_000 byte 2 was rd_b4_wr
  //(cp_log_000_rst_val_chk): Cover that DEV_CAR_OVRD is non-default and log_000 was rd_b4_wr
  //(cp_log_004_rd_b4_wr): Cover that each byte of log_004 was read before it was written
  //(cp_log_004_rd_aftr_wr): Cover that each byte of log_004 was read after it was written
  //(cp_log_004_rst_val_chk): Cover that DEV_CAR_OVRD is non-default and log_004 was rd_b4_wr
  //(cp_log_008_rd_b4_wr): Cover that each byte of log_008 was read before it was written
  //(cp_log_008_rd_aftr_wr): Cover that each byte of log_008 was read after it was written
  //(cp_log_008_3_rst_val_chk): Cover that ASSY_ID is non-default and log_008 byte 3 was rd_b4_wr
  //(cp_log_008_2_rst_val_chk): Cover that ASSY_ID is non-default and log_008 byte 2 was rd_b4_wr
  //(cp_log_008_1_rst_val_chk): Cover that ASSY_VENDOR is non-default and log_008 byte 3 was rd_b4_wr
  //(cp_log_008_0_rst_val_chk): Cover that ASSY_VENDOR is non-default and log_008 byte 2 was rd_b4_wr
  //(cp_log_00c_rd_b4_wr): Cover that each byte of log_00c was read before it was written
  //(cp_log_00c_rd_aftr_wr): Cover that each byte of log_00c was read after it was written
  //(cp_log_00c_3_rst_val_chk): Cover that ASSY_REV is non-default and log_00c byte 3 was rd_b4_wr
  //(cp_log_00c_2_rst_val_chk): Cover that ASSY_REV is non-default and log_00c byte 2 was rd_b4_wr
  //(cp_log_00c_1_rst_val_chk): Cover that PHY_EF_PTR is non-default and log_00c byte 3 was rd_b4_wr
  //(cp_log_00c_0_rst_val_chk): Cover that PHY_EF_PTR is non-default and log_00c byte 2 was rd_b4_wr
  //(cp_log_010_rd_b4_wr): Cover that each byte of log_010 was read before it was written
  //(cp_log_010_rd_aftr_wr): Cover that each byte of log_010 was read after it was written
  //(cp_log_010_bit31_rst_val_chk): Cover that PE_BRIDGE is non-default and log_010 bit 31 was rd_b4_wr
  //(cp_log_010_bit30_rst_val_chk): Cover that PE_MEMORY is non-default and log_010 bit 30 was rd_b4_wr
  //(cp_log_010_bit29_rst_val_chk): Cover that PE_PROC is non-default and log_010 bit 29 was rd_b4_wr
  //(cp_log_010_bit28_rst_val_chk): Cover that PE_SWITCH is non-default and log_010 bit 28 was rd_b4_wr
  //(cp_log_010_bit5_rst_val_chk): Cover that CRF_SUPPORT is non-default and log_010 bit 5 was rd_b4_wr
  //(cp_log_010_bit4_rst_val_chk): Cover that DEVICEID_WIDTH is non-default and log_010 bit 4 was rd_b4_wr
  //(cp_log_018_rd_b4_wr): Cover that each byte of log_018 was read before it was written
  //(cp_log_018_rd_aftr_wr): Cover that each byte of log_018 was read after it was written
  //(cp_log_018_bit15_rst_val_chk): Cover that INIT_NREAD is non-default and log_018 bit 15 was rd_b4_wr
  //(cp_log_018_bit14_rst_val_chk): Cover that INIT_NWRITE is non-default and log_018 bit 14 was rd_b4_wr
  //(cp_log_018_bit13_rst_val_chk): Cover that INIT_SWRITE is non-default and log_018 bit 13 was rd_b4_wr
  //(cp_log_018_bit12_rst_val_chk): Cover that INIT_NWRITE_R is non-default and log_018 bit 12 was rd_b4_wr
  //(cp_log_018_bit11_rst_val_chk): Cover that INIT_MSG is non-default and log_018 bit 11 was rd_b4_wr
  //(cp_log_018_bit10_rst_val_chk): Cover that INIT_DB is non-default and log_018 bit 10 was rd_b4_wr
  //(cp_log_018_1_rst_val_chk): Cover that INIT_ATOMIC is non-default and log_018 byte 1 was rd_b4_wr
  //(cp_log_018_0_rst_val_chk): Cover that INIT_ATOMIC is non-default and log_018 byte 0 was rd_b4_wr
  //(cp_log_01c_rd_b4_wr): Cover that each byte of log_01c was read before it was written
  //(cp_log_01c_rd_aftr_wr): Cover that each byte of log_01c was read after it was written
  //(cp_log_01c_bit15_rst_val_chk): Cover that TARGET_NREAD is non-default and log_01c bit 15 was rd_b4_wr
  //(cp_log_01c_bit14_rst_val_chk): Cover that TARGET_NWRITE is non-default and log_01c bit 14 was rd_b4_wr
  //(cp_log_01c_bit13_rst_val_chk): Cover that TARGET_SWRITE is non-default and log_01c bit 13 was rd_b4_wr
  //(cp_log_01c_bit12_rst_val_chk): Cover that TARGET_NWRITE_R is non-default and log_01c bit 12 was rd_b4_wr
  //(cp_log_01c_bit11_rst_val_chk): Cover that TARGET_MSG is non-default and log_01c bit 11 was rd_b4_wr
  //(cp_log_01c_bit10_rst_val_chk): Cover that TARGET_DB is non-default and log_01c bit 10 was rd_b4_wr
  //(cp_log_01c_1_rst_val_chk): Cover that TARGET_ATOMIC is non-default and log_01c byte 1 was rd_b4_wr
  //(cp_log_01c_0_rst_val_chk): Cover that TARGET_ATOMIC is non-default and log_01c byte 0 was rd_b4_wr
  //(cp_log_04c_rd_b4_wr): Cover that each byte of log_04c was read before it was written
  //(cp_log_04c_rd_aftr_wr): Cover that each byte of log_04c was read after it was written
  //(cp_log_058_rd_b4_wr): Cover that each byte of log_058 was read before it was written
  //(cp_log_058_rd_aftr_wr): Cover that each byte of log_058 was read after it was written
  //(cp_log_05c_rd_b4_wr): Cover that each byte of log_05c was read before it was written
  //(cp_log_05c_rd_aftr_wr): Cover that each byte of log_05c was read after it was written
  //(cp_log_05c_3_rst_val_chk): Cover that LCSBA is non-default and log_05c byte 3 was rd_b4_wr
  //(cp_log_05c_3_rst_val_chk_no_lcsba): Cover that LCSBA_SUPPORT is non-default and log_05c byte 3 was rd_b4_wr
  //(cp_log_05c_2_rst_val_chk): Cover that LCSBA is non-default and log_05c byte 2 was rd_b4_wr
  //(cp_log_05c_2_rst_val_chk_no_lcsba): Cover that LCSBA_SUPPORT is non-default and log_05c byte 3 was rd_b4_wr
  //(cp_log_060_rd_b4_wr): Cover that each byte of log_060 was read before it was written
  //(cp_log_060_rd_aftr_wr): Cover that each byte of log_060 was read after it was written
  //(cp_log_060_2_rst_val_chk): Cover that DEVICEID is non-default and log_060 byte 2 was rd_b4_wr
  //(cp_log_060_1_rst_val_chk): Cover that DEVICEID is non-default and log_060 byte 1 was rd_b4_wr
  //(cp_log_060_0_rst_val_chk): Cover that DEVICEID is non-default and log_060 byte 0 was rd_b4_wr
  //(cp_log_068_rd_b4_wr): Cover that each byte of log_068 was read before it was written
  //(cp_log_068_rd_aftr_wr): Cover that each byte of log_068 was read after it was written
  //(cp_log_06c_rd_b4_wr): Cover that each byte of log_06c was read before it was written
  //(cp_log_06c_rd_aftr_wr): Cover that each byte of log_06c was read after it was written

  // Register read data when address is safe
  // No reset needed since data is not sampled until valid
  always @(posedge log_clk) begin
    if (CCA_sync_re) begin
      case (CCA_cfg_raddr[15:0])
        LOG_000    : LCR_core_rdata <= #TCQ csr_log_000;
        LOG_004    : LCR_core_rdata <= #TCQ csr_log_004;
        LOG_008    : LCR_core_rdata <= #TCQ csr_log_008;
        LOG_00C    : LCR_core_rdata <= #TCQ csr_log_00c;
        LOG_010    : LCR_core_rdata <= #TCQ csr_log_010;
        LOG_014    : LCR_core_rdata <= #TCQ csr_log_014;
        LOG_018    : LCR_core_rdata <= #TCQ csr_log_018;
        LOG_01C    : LCR_core_rdata <= #TCQ csr_log_01c;
        LOG_04C    : LCR_core_rdata <= #TCQ csr_log_04c;
        LOG_058    : LCR_core_rdata <= #TCQ csr_log_058;
        LOG_05C    : LCR_core_rdata <= #TCQ csr_log_05c;
        LOG_060    : LCR_core_rdata <= #TCQ csr_log_060;
        LOG_068    : LCR_core_rdata <= #TCQ csr_log_068;
        LOG_06C    : LCR_core_rdata <= #TCQ csr_log_06c;
        // Return data of all 0's if read to unimplemented space
        default    : LCR_core_rdata <= #TCQ 32'b0;
      endcase
    end
  end

  // }}} End Read Data Assembly ------------


endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/log/log_cfg/srio_gen2_v4_1_16_log_cfg_top.v#3 $
//----------------------------------------------------------------------
//
// LOG_CFG
// Description:
// This module contains the configuration registers for the LOG layer.
//
// It uses an AXI-Lite interface to the Configuration Fabric, and has a
// core interface for transfer of control and status information.
//
// No clock relationship between cfg_clk and the log_clk is assumed.
//
// Hierarchy:
// LOG_TOP
//  |______LOG_CFG_TOP <-- this module
//            |______CFG_AXI (in hdl/common/)
//            |______LOG_CFG_REG
// ---------------------------------------------------------------------
`timescale 1ps/1ps

// ------------------------------------------------
// below attribute is added to supress the synthesis warnings in vivado tool 8:3332
(* DowngradeIPIdentifiedWarnings="yes" *)
// ------------------------------------------------

module srio_gen2_v4_1_16_log_cfg_top
  #(
      parameter TCQ   = 100,
      parameter HW_ARCH         = 2,          // Device {V5LXT(0), V5FXT(1), V6LXT(2), V6CXT(3), S6LXT(4)}
      parameter DEVICEID_WIDTH  = 8,          // Source/Destination ID width {8,16}
      parameter DEVICEID        = 16'h00FF,   // Reset value for Device ID {16'h0000-16'hFFFF}
      parameter INIT_NREAD      = 1,          // Core may initiate NREAD transactions {0,1}
      parameter INIT_NWRITE     = 1,          // Core may initiate NWRITE transactions {0,1}
      parameter INIT_SWRITE     = 1,          // Core may initiate SWRITE transactions {0,1}
      parameter INIT_NWRITE_R   = 1,          // Core may initiate NWRITE_R transactions {0,1}
      parameter INIT_DB         = 1,          // Core may initiate Doorbell transactions {0,1}
      parameter INIT_DS         = 1,          // Core may initiate Data-Streaming transactions {0,1}
      parameter INIT_ATOMIC     = 1,          // Core may initiate ATOMIC transactions {0,1}
      parameter MSG_INIT_SINGLE = 1,          // Core may initiate single-segment message transactions {0,1}
      parameter MSG_INIT_MULTI  = 1,          // Core may initiate multiple-segment message transactions {0,1}
      parameter TARGET_NREAD    = 1,          // Core may sink NREAD transactions {0,1}
      parameter TARGET_NWRITE   = 1,          // Core may sink NWRITE transactions {0,1}
      parameter TARGET_SWRITE   = 1,          // Core may sink SWRITE transactions {0,1}
      parameter TARGET_NWRITE_R = 1,          // Core may sink NWRITE_R transactions {0,1}
      parameter TARGET_DB       = 1,          // Core may sink Doorbell transactions {0,1}
      parameter TARGET_DS       = 1,          // Core may initiate Data-Streaming transactions {0,1}
      parameter TARGET_ATOMIC   = 1,          // Core may sink ATOMIC transactions {0,1}
      parameter MSG_SINK_SINGLE = 1,          // Core may sink single-segment message transactions {0,1}
      parameter MSG_SINK_MULTI  = 1,          // Core may sink multiple-segment message transactions {0,1}
      parameter CRF_SUPPORT     = 1,          // If set, the core supports use of the CRF flag {0,1}
      parameter DEVID_CAR       = 32'h00000000,   // Reset value for Device Identity CAR {32�h00000000�?32�hFFFFFFFF}
      parameter DEVINFO_CAR     = 32'h00000000,   // Reset value for Device Info CAR {32�h00000000�?32�hFFFFFFFF}
      parameter DEV_CAR_OVRD    = 0,              // If 1, DEV*CAR param values used {0,1}
      parameter LCSBA_SUPPORT   = 1,          // If set, I/O transactions can be rerouted to the maint port {0,1}
      parameter LCSBA           = 10'h3FF,    // Reset value for LCSBA register {10'h0-10'h3FF}
      parameter ASSY_ID         = 16'h0000,   // Assembly ID from GUI {16'h0000-16'hFFFF}
      parameter ASSY_VENDOR     = 16'h0000,   // Assembly Vendor ID from GUI {16'h0000-16'hFFFF}
      parameter ASSY_REV        = 16'h0000,   // Assembly Revision from GUI {16'h0000-16'hFFFF}
      parameter PE_BRIDGE       = 0,          // Processing Element contains Bridge functionality {0,1}
      parameter PE_MEMORY       = 1,          // Processing Element contains Memory functionality {0,1}
      parameter PE_PROC         = 0,          // Processing Element contains Processor functionality {0,1}
      parameter PE_SWITCH       = 0,          // Processing Element contains Switch functionality {0,1}
      parameter PHY_EF_PTR      = 16'h0100  // Location of PHY ext features {0x0100+}
  )(
    // {{{ Port Declarations ---------------
    // System Signals
    input             log_clk,                // LOG interface clock
    input             log_rst,                // Reset for LOG clock Domain
    input             cfg_clk,                // CFG Interface user clock
    input             cfg_rst,                // Reset for CFG clk domain

    // User Interface
    output     [15:0] LC_deviceid,            // Current Device ID - Used as SourceID for transmitted transactions

    // LOG Arb Interface
    output     [9:0]  LC_lcsba,               // Local Configuration Base Address register mask value

    // Configuration Fabric Interface
    input             CF_cfgl_awvalid,        // Write Address Valid
    output            LC_cfgl_awready,        // Write Address Port Ready
    input      [23:0] CF_cfgl_awaddr,         // Write Address
    input             CF_cfgl_wvalid,         // Write Data Valid
    output            LC_cfgl_wready,         // Write Data Port Ready
    input      [31:0] CF_cfgl_wdata,          // Write Data
    input      [3:0]  CF_cfgl_wstrb,          // Write Data Byte Enables
    output            LC_cfgl_bvalid,         // Write Response Valid
    input             CF_cfgl_bready,         // Write Response Fabric Ready
    input             CF_cfgl_arvalid,        // Read Address Valid
    output            LC_cfgl_arready,        // Read Address Port Ready
    input      [23:0] CF_cfgl_araddr,         // Read Address
    output            LC_cfgl_rvalid,         // Read Response Valid
    input             CF_cfgl_rready,         // Read Response Fabric Ready
    output     [31:0] LC_cfgl_rdata           // Read Data
    // }}} End Port Declarations -----------
  );

  // {{{ Wire Declarations -----------------
  wire              CCA_sync_cfg_rst;         // cfg_rst sync'ed to log_clk
  wire       [23:0] CCA_cfg_waddr;            // Write Address
  wire       [31:0] CCA_cfg_wdata;            // Write Data
  wire       [3:0]  CCA_cfg_wstrb;            // Write Data Byte Enables
  wire              CCA_sync_we;              // Synchronized write enable
  wire       [23:0] CCA_cfg_raddr;            // Read Address
  wire              CCA_sync_re;              // Synchronized Read Enable
  wire       [31:0] LCR_core_rdata;           // Read Data
  // }}} End Wire Declarations -------------


  // {{{ log_cfg_axi inst ------------------
  // Instantiate the generic cfg interface, which contains the clock domain
  // crossing from cfg_clk to log_clk, as well as the AXI-Lite interface to
  // the CFG Fabric
  srio_gen2_v4_1_16_cfg_axi
    #(
      .TCQ                       (TCQ))
    log_cfg_axi_inst
     (.core_clk                  (log_clk),
      .cfg_clk                   (cfg_clk),
      .cfg_rst                   (cfg_rst),
      .CF_awvalid                (CF_cfgl_awvalid),
      .CCA_awready               (LC_cfgl_awready),
      .CF_awaddr                 (CF_cfgl_awaddr),
      .CF_wvalid                 (CF_cfgl_wvalid),
      .CCA_wready                (LC_cfgl_wready),
      .CF_wdata                  (CF_cfgl_wdata),
      .CF_wstrb                  (CF_cfgl_wstrb),
      .CCA_bvalid                (LC_cfgl_bvalid),
      .CF_bready                 (CF_cfgl_bready),
      .CF_arvalid                (CF_cfgl_arvalid),
      .CCA_arready               (LC_cfgl_arready),
      .CF_araddr                 (CF_cfgl_araddr),
      .CCA_rvalid                (LC_cfgl_rvalid),
      .CF_rready                 (CF_cfgl_rready),
      .CCA_rdata                 (LC_cfgl_rdata),
      .CCA_sync_cfg_rst          (CCA_sync_cfg_rst),
      .CCA_cfg_waddr             (CCA_cfg_waddr),
      .CCA_cfg_wdata             (CCA_cfg_wdata),
      .CCA_cfg_wstrb             (CCA_cfg_wstrb),
      .CCA_sync_we               (CCA_sync_we),
      .CCA_cfg_raddr             (CCA_cfg_raddr),
      .CCA_sync_re               (CCA_sync_re),
      .CC_core_rdata             (LCR_core_rdata));
  // }}} End log_cfg_axi inst --------------

  // {{{ log_cfg_reg inst ------------------
  //----------------------------------------
  srio_gen2_v4_1_16_log_cfg_reg
    #(.TCQ                       (TCQ),
      .HW_ARCH                   (HW_ARCH),
      .DEVICEID_WIDTH            (DEVICEID_WIDTH),
      .DEVICEID                  (DEVICEID),
      .INIT_NREAD                (INIT_NREAD),
      .INIT_NWRITE               (INIT_NWRITE),
      .INIT_SWRITE               (INIT_SWRITE),
      .INIT_NWRITE_R             (INIT_NWRITE_R),
      .INIT_DB                   (INIT_DB),
      .INIT_DS                   (INIT_DS),
      .INIT_ATOMIC               (INIT_ATOMIC),
      .MSG_INIT_SINGLE           (MSG_INIT_SINGLE),
      .MSG_INIT_MULTI            (MSG_INIT_MULTI),
      .CRF_SUPPORT               (CRF_SUPPORT),
      .TARGET_NREAD              (TARGET_NREAD),
      .TARGET_NWRITE             (TARGET_NWRITE),
      .TARGET_SWRITE             (TARGET_SWRITE),
      .TARGET_NWRITE_R           (TARGET_NWRITE_R),
      .TARGET_DB                 (TARGET_DB),
      .TARGET_DS                 (TARGET_DS),
      .TARGET_ATOMIC             (TARGET_ATOMIC),
      .MSG_SINK_SINGLE           (MSG_SINK_SINGLE),
      .MSG_SINK_MULTI            (MSG_SINK_MULTI),
      .DEVID_CAR                 (DEVID_CAR),
      .DEVINFO_CAR               (DEVINFO_CAR),
      .DEV_CAR_OVRD              (DEV_CAR_OVRD),
      .LCSBA_SUPPORT             (LCSBA_SUPPORT),
      .LCSBA                     (LCSBA),
      .ASSY_ID                   (ASSY_ID),
      .ASSY_VENDOR               (ASSY_VENDOR),
      .ASSY_REV                  (ASSY_REV),
      .PE_BRIDGE                 (PE_BRIDGE),
      .PE_MEMORY                 (PE_MEMORY),
      .PE_PROC                   (PE_PROC),
      .PE_SWITCH                 (PE_SWITCH),
      .PHY_EF_PTR                (PHY_EF_PTR))
    log_cfg_reg_inst
     (.log_clk                   (log_clk),
      .log_rst                   (log_rst),
      .CCA_sync_cfg_rst          (CCA_sync_cfg_rst),
      .LCR_lcsba                 (LC_lcsba),
      .LCR_deviceid              (LC_deviceid),
      .CCA_cfg_waddr             (CCA_cfg_waddr),
      .CCA_cfg_wdata             (CCA_cfg_wdata),
      .CCA_cfg_wstrb             (CCA_cfg_wstrb),
      .CCA_sync_we               (CCA_sync_we),
      .CCA_cfg_raddr             (CCA_cfg_raddr),
      .CCA_sync_re               (CCA_sync_re),
      .LCR_core_rdata            (LCR_core_rdata));
  // }}} End log_cfg_reg inst

endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}


//----------------------------------------------------------------------
// $Id: //IP3/DEV/hw/srio_gen2/srio_gen2_v4_1_16/hdl/log/log_maint/srio_gen2_v4_1_16_log_maint.v#1 $
//----------------------------------------------------------------------
//
// LOG_MAINT
// Description:
// This module accepts maintenance requests from the user and the link
// partner, routes them to the Configuration Fabric or to the Arbiter
// for transmission on the link, and returns the response.
//
// Hierarchy:
// LOG_TOP
//    |___LOG_MAINT
// ---------------------------------------------------------------------

`timescale 1ps/1ps

module srio_gen2_v4_1_16_log_maint
#(parameter TCQ                  =      100,  // in ps
  parameter DEVICEID_WIDTH       =        8,  // Indicates Source/Dest ID width {8, 16}
  parameter TARGET_NREAD         =        1,  // If 1, core may sink NRead transactions {0, 1}
  parameter TARGET_NWRITE        =        1,  // If 1, core may sink NWrite transactions {0, 1}
  parameter TARGET_NWRITE_R      =        1,  // If 1, core may sink NWrite_R transactions {0, 1}
  parameter CRF_SUPPORT          =        1,  // If set, the core supports use of the CRF flag {0,1}
  parameter MAINT_SOURCE         =        1,  // If 1, core may source maintenance transactions {0, 1}
  parameter LCSBA_SUPPORT        =        1,  // If 1, indicates the LCSBA is used {0, 1}
  parameter VC                   =        0)  // If 1, VC is supported
(
  // {{{ port declarations -----------------
  // System Interface
  input                 log_clk,              // LOG interface clock
  input                 log_rst,              // Reset for LOG clock Domain
  input                 maintr_rst,           // Reset for maintr interface, on LOG clock Domain

  // LOG User Maintenance Interface
  // AXI-Lite Slave
  //----------------------------------------
  // Write Address Channel
  input                 UG_maintr_awvalid,    // Write Address Valid
  output reg            LR_maintr_awready,    // Ready for Write Address
  input      [31:0]     UG_maintr_awaddr,     // Write Address

  // Write Data Channel
  input                 UG_maintr_wvalid,     // Write Data Valid
  output reg            LR_maintr_wready,     // Ready for Write Data
  input      [31:0]     UG_maintr_wdata,      // Write Data

  // Write Response Channel
  output reg            LR_maintr_bvalid,     // Write Response Valid
  input                 UG_maintr_bready,     // Write Response Fabric Ready
  output reg [1:0]      LR_maintr_bresp = 0,  // Write Response

  // Read Address Channel
  input                 UG_maintr_arvalid,    // Read Command Valid
  output reg            LR_maintr_arready,    // Read Port Ready
  input      [31:0]     UG_maintr_araddr,     // Read Address

  // Read Response Channel
  output reg            LR_maintr_rvalid,     // Read Response Valid
  input                 UG_maintr_rready,     // Read Response Fabric Ready
  output reg [31:0]     LR_maintr_rdata = 0,  // Read Data
  output reg [1:0]      LR_maintr_rresp = 0,  // Read Response

  // Maintenace/Config Fabric Interface
  // AXI-Lite Master
  //----------------------------------------
  // Write Address Channel
  output reg            LR_cfgr_awvalid,      // Write Address Valid
  input                 CF_cfgr_awready,      // Ready for Write Address
  output reg [23:0]     LR_cfgr_awaddr,       // Write Address
  output     [2:0]      LR_cfgr_awprot,       // Write Protection (Tied to 0)

  // Write Data Channel
  output reg            LR_cfgr_wvalid,       // Write Data Valid
  input                 CF_cfgr_wready,       // Ready for Write Data
  output reg [31:0]     LR_cfgr_wdata,        // Write Data
  output     [3:0]      LR_cfgr_wstrb,        // Write Data byte enables

  // Write Response Channel
  input                 CF_cfgr_bvalid,       // Write Response Valid
  output reg            LR_cfgr_bready,       // Write Response Fabric Ready
  input      [1:0]      CF_cfgr_bresp,        // Write Response

  // Read Address Channel
  output reg            LR_cfgr_arvalid,      // Read Command Valid
  input                 CF_cfgr_arready,      // Read Port Ready
  output reg [23:0]     LR_cfgr_araddr,       // Read Address
  output     [2:0]      LR_cfgr_arprot,       // Read Protection (Tied to 0)

  // Read Response Channel
  input                 CF_cfgr_rvalid,       // Read Response Valid
  output reg            LR_cfgr_rready,       // Read Response Fabric Ready
  input      [31:0]     CF_cfgr_rdata,        // Read Data
  input      [1:0]      CF_cfgr_rresp,        // Read Response

  // LOG Arb TX Request Interface
  // AXI-Streaming Master
  //----------------------------------------
  output reg            LR_lrtx_req_tvalid=0, // Valid packet beat
  input                 LA_lrtx_req_tready,   // Packet beat accepted
  output reg [63:0]     LR_lrtx_req_tdata,    // Packet data
  output     [7:0]      LR_lrtx_req_tkeep,    // Valid bytes in this beat, only valid on last
  output reg            LR_lrtx_req_tlast=0,  // Last beat
  output reg [39:0]     LR_lrtx_req_tuser,    // {SrcID, DestID, 2'b0, HELLO_FMT (1), Response (0), 1'b0, CRF, 1'b0}

  // LOG Arb TX Response Interface
  // AXI-Streaming Master
  //----------------------------------------
  output reg            LR_lrtx_resp_tvalid=0,// Valid packet beat
  input                 LA_lrtx_resp_tready,  // Packet beat accepted
  output reg [63:0]     LR_lrtx_resp_tdata,   // Packet data
  output     [7:0]      LR_lrtx_resp_tkeep,   // Valid bytes in this beat, only valid on last
  output reg            LR_lrtx_resp_tlast=0, // Last beat
  output reg [39:0]     LR_lrtx_resp_tuser,   // {SrcID, DestID, 2'b0, HELLO_FMT (1), Response (1), 1'b0, CRF, 1'b0}

  // LOG Arb RX Interface
  // AXI-Streaming Slave
  //----------------------------------------
  input                 LA_lrrx_tvalid,       // Valid packet beat
  output reg            LR_lrrx_tready,       // Packet beat accepted
  input      [63:0]     LA_lrrx_tdata,        // Packet data
  input      [7:0]      LA_lrrx_tkeep,        // Valid bytes in this beat, only valid on last
  input                 LA_lrrx_tlast,        // Last beat
  input      [39:0]     LA_lrrx_tuser,        // {SrcID, DestID, 2'b0, HELLO_FMT (1), Response, 1'b0, CRF, 1'b0}

  // LOG CFG Interface
  //----------------------------------------
  input      [15:0]     LC_deviceid           // Device ID from Device Identity CSR to be used as srcID
  );
  // }}} end port declarations -------------

  // {{{ Local Parameters
  // Spec defined parameters
  // ------------------------------------------------------------
  // Ftype
  localparam FTYPE_NREAD    = 4'b0010;
  localparam FTYPE_NWRITE   = 4'b0101;
  localparam FTYPE_SWRITE   = 4'b0110;
  localparam FTYPE_MAINT    = 4'b1000;
  localparam FTYPE_RESP     = 4'b1101;
  // Ttype
  localparam TTYPE_NREAD    = 4'b0100;
  localparam TTYPE_NWRITE   = 4'b0100;
  localparam TTYPE_NWRITE_R = 4'b0101;
  localparam TTYPE_MREQR    = 4'b0000;
  localparam TTYPE_MREQW    = 4'b0001;
  localparam TTYPE_MRESPR   = 4'b0010;
  localparam TTYPE_MRESPW   = 4'b0011;
  localparam TTYPE_RESPW    = 4'b0000;
  localparam TTYPE_RESPR    = 4'b1000;
  // Status
  localparam STAT_DONE      = 4'b0000;
  localparam STAT_ERR       = 4'b0111;
  // TT
  localparam TT             = (DEVICEID_WIDTH == 8) ? 2'b0 : 2'b01; // tt field
  // Encodings for sending signals
  localparam SENDING_NONE   = 2'b00;
  localparam SENDING_READ   = 2'b01;
  localparam SENDING_WRITE  = 2'b10;
  // Offset of Maintenance Request Information CSR
  localparam CSR_INFO_REG   = 24'h01_0100; // Offset 0x100 within Implementation-Defined space
  // }}} end Local Parameters

  // {{{ Wire Declarations
  reg                       log_rst_q  = 1;     // Registered version of log_rst
  reg                       maintrlog_rst_q = 1;// Registered log_rst || maintr_rst, clears outstanding maintr request
  reg                       maintrlog_rst_qq= 1;// Registered maintrlog_rst_q, re-sets readys after reset
  // Signals for User Interface
  wire                      lru_aractive;       // User Read Address channel active (ready && valid)
  reg                       lru_aractive_q;     // Registered version of lru_aractive
  wire                      lru_ractive;        // User Read Response channel active (ready && valid)
  reg  [31:0]               lru_raddr;          // User read address
  wire                      lru_awactive;       // User Write Address channel active (ready && valid)
  wire                      lru_wactive;        // User Write Data channel active (ready && valid)
  wire                      lru_bactive;        // User Write Response channel active (ready && valid)
  reg  [31:0]               lru_waddr;          // User write address
  reg  [31:0]               lru_wdata;          // User write data
  reg                       lru_got_waddr;      // A User write address has been accepted
  reg                       lru_got_wdata;      // User write data had been accepted
  // Signals for Arbiter RX Interface
  wire                      lrr_active;         // lrrx interface active (ready && valid)
  reg                       lrr_tlast_hold;     // LA_lrrx_tlast registered on lrr_active
  reg                       lrr_sof_hold;       // Registered version of lrr_sof
  wire                      lrr_sof;            // First DWORD of packet accepted from arbiter
  wire                      lrr_last;           // Last DWORD of packet accepted from arbiter
  wire [7:0]                lrr_tid;            // Received TID
  wire [3:0]                lrr_ftype;          // FTYPE of packet on lrrx interface
  wire [3:0]                lrr_ttype;          // TTYPE of packet on lrrx interface
  wire [1:0]                lrr_prio;           // The priority field of a received packet
  wire                      lrr_crf;            // The CRF for a received packet
  wire [7:0]                lrr_size;           // The size of a received packet
  wire                      lrr_ok;             // Status of received Response
  wire [23:0]               lrr_addr;           // The address from the received packet
  reg                       lrr_ok_hold;        // Registered version of status of received Response
  reg                       lrr_addr_hold;      // Registered version of address from the received packet
  wire                      lrr_read;           // Transaction on lrrx interface is a read request
  wire                      lrr_write;          // Transaction on lrrx interface is a write request
  wire                      lrr_rresp;          // Transaction on lrrx interface is a read response
  wire                      lrr_wresp;          // Transaction on lrrx interface is a write response
  wire                      lrr_req_sof;        // First DWORD of a request packet accepted from arbiter
  reg                       lrr_req_pending;    // A request from the arb is pending
  wire                      lrr_set_rdy;        // Used to set the lrrx_ready signal
  // Signals for Config Fabric Interface
  wire                      lrc_aractive;       // Config Fabric Read Address channel active (ready && valid)
  wire                      lrc_ractive;        // Config Fabric Read Response channel active (ready && valid)
  reg  [31:0]               lrc_rdata;          // Config Fabrid read data
  reg  [1:0]                lrc_rresp;          // Config Fabric read response
  reg                       lrc_got_rresp;      // A read response has been received from the Config Fabric
  wire                      lrc_awactive;       // Config Fabric Write Address channel active (ready && valid)
  wire                      lrc_wactive;        // Config Fabric Write Data channel active (ready && valid)
  wire                      lrc_bactive;        // Config Fabric Write Response channel active (ready && valid)
  reg  [1:0]                lrc_wresp;          // Config Fabric write response
  reg                       lrc_got_wresp;      // A write response has been received from the Config Fabric
  // Signals for Request Info Register
  reg                       lri_req_vc;         // The VC field for outgoing requests, from Req Info reg
  reg  [1:0]                lri_req_prio;       // The prio field for outgoing requests, from Req Info reg
  reg                       lri_req_crf;        // The CRF field for outgoing requests, from Req Info reg
  reg  [15:0]               lri_req_destid;     // The Destination ID field for outgoing requests, from Req Info reg
  reg  [7:0]                lri_req_next_tid;   // The TID field for outgoing requests (increments from base_tid)
  wire [31:0]               lri_csr_lr_000;     // The value of the Request Info reg for register reads
  // Signals for User Read Manager
  wire                      lrm_ur_info;        // The user read targets the LOG Request Info Register
  wire                      lrm_ur_local;       // The read transaction from the user targets the local config space
  wire                      lrm_ur_remote;      // The read transaction from the user targets the remote config space
  reg                       lrm_ur_info_pend;   // The pending user read targets the LOG Request Info Register
  reg                       lrm_ur_local_pend;  // The pending read transaction from the user targets the local config space
  reg                       lrm_ur_remote_pend; // The pending read transaction from the user targets the remote config space
  reg                       lrm_ur_read_lock;   // The user "owns" the read channels of the Config Fabric interface
  reg                       lrm_ur_read_lock_q; // Registered version of lrm_ur_read_lock
  wire                      lrm_ur_read_cfg;    // A user CF read is ready
  reg                       lrm_ur_rreq_gen;    // The user read manager is requesting a read MREQ to be transmitted
  wire [7:0]                lrm_ur_hopcount;    // Hopcount for user read (decrement MSB of user address)
  reg  [7:0]                lrm_ur_tid;         // TID assigned to user read (based on Req Info register)
  reg                       lrm_ur_tid_match;   // Identifies a match of the TID of the received response with the req
  wire                      lrm_ur_got_rresp;   // A read response for the user is available
  wire [1:0]                lrm_ur_rresp;       // Read response for the user
  wire [31:0]               lrm_ur_rdata;       // Read data (as part of read response) for the user
  // Signals for User Write Manager
  wire                      lrm_uw_info;        // The user write targets the LOG Request Info Register
  wire                      lrm_uw_local;       // The write transaction from the user targets the local config space
  wire                      lrm_uw_remote;      // The write transaction from the user targets the remote config space
  reg                       lrm_uw_info_pend;   // A user write targeting the LOG Request Info Register is pending
  reg                       lrm_uw_local_pend;  // A user write targeting the local config space is pending
  reg                       lrm_uw_remote_pend; // A user write targeting the remote config space is pending
  reg                       lrm_uw_write_lock;  // The User Write Manager "owns" the write channels of the CF interface
  reg                       lrm_uw_write_lock_q;// Registered version of lrm_ur_write_lock
  wire                      lrm_uw_write_cfg;   // A user CF write is ready
  reg                       lrm_uw_info_reg_wen;// Write enable for Request Info register
  reg                       lrm_uw_wreq_gen;    // The user write manager is requesting a write MREQ to be transmitted
  reg  [7:0]                lrm_uw_tid;         // TID assigned to user write (based on Req Info register)
  wire [7:0]                lrm_uw_hopcount;    // Hopcount for user write (decrement MSB of user address)
  reg                       lrm_uw_tid_match;   // Identifies a match of the TID of the received response with the req
  wire                      lrm_uw_got_wresp;   // A write response for the user is available
  wire [1:0]                lrm_uw_wresp;       // Write response for the user
  // Signals for External Request Manager
  reg                       lrm_ext_read_lock;  // The External Request Manager "owns" the read CF interface
  reg                       lrm_ext_write_lock; // The External Request Manager "owns" the write CF interface
  wire                      lrm_ext_read_rdy;   // An external read is ready (last write beat accepted from arb)
  wire                      lrm_ext_write_rdy;  // An external write is ready (last write beat accepted from arb)
  wire                      lrm_ext_size_ok;    // The external request's size is valid
  wire                      lrm_ext_type_ok;    // The external request's TTYPE is valid
  wire                      lrm_ext_req_ok;     // The external request is valid
  reg                       lrm_ext_req_ok_hold;// lrm_ext_req_ok captured on sof for use after sof
  reg                       lrm_ext_no_resp;    // The external request does not require a response
  wire                      lrm_ext_info_reg_ren;   // Read enable for Request Info register
  wire                      lrm_ext_read_cfg;   // An external CF read is ready
  wire                      lrm_ext_read_err;   // The size or TTYPE of the external request is invalid
  reg                       lrm_ext_info_read;  // The external read targets the Req Info reg
  wire                      lrm_ext_got_waddr;  // Flag used to overwrite the addr to the CF on beat 2
  reg                       lrm_ext_info_reg_write; // The write on lrr targets the maint request info register
  wire                      lrm_ext_info_reg_wen;   // Write enable for Request Info register
  wire                      lrm_ext_write_cfg;  // An external write is ready for the CF interface
  wire                      lrm_ext_write_err;  // The external write request has an error
  wire                      lrm_ext_cfg_rresp;  // A read response is available from the Config Fabric
  wire                      lrm_ext_cfg_wresp;  // A write response is available from the Config Fabric
  reg  [3:0]                lrm_ext_resp_ftype; // The FTYPE for the response to the external request
  reg  [3:0]                lrm_ext_resp_ttype; // The TTYPE for the response to the external request
  wire [1:0]                lrm_ext_resp_prio;  // The priority for the response to the external request
  reg                       lrm_ext_resp_err;   // The status for the response to the external request
  reg                       lrm_ext_rresp_gen;  // Generate a read response packet for transmit
  reg                       lrm_ext_wresp_gen;  // Generate a write response packet for transmit
  // Signals for Response Generator
  wire                      lrs_valid;          // The response generator signals (e.g. lrs_pkt) are valid
  wire                      lrs_resp_w_data;    // The response has data (i.e. unerrored read response)
  wire                      lrs_header_stage;   // Generating the header for a response
  reg                       lrs_data_stage;     // Generating the data for a response
  wire                      lrs_active;         // The lrtx_resp interface is active (ready && valid)
  wire                      lrs_resp_sent;      // A response was accepted for transmission by the arb
  // Signals for Request Generator
  wire                      lrq_valid;          // A request is in progress
  wire                      lrq_start;          // The request generator is creating a new request
  wire [1:0]                lrq_pktsel;         // The packet type to generate
  reg  [1:0]                lrq_pktsel_hold;    // lrq_pktsel registered on the first beat
  wire [1:0]                lrq_sending;        // The packet type being generated
  wire [3:0]                lrq_ttype;          // The request TTYPE
  wire [7:0]                lrq_size;           // The request size
  wire [7:0]                lrq_hopcount;       // The request hopcount
  wire [23:0]               lrq_addr;           // The request address
  wire [63:0]               lrq_header;         // The header selected based on request type
  wire [63:0]               lrq_data;           // The data for a write request
  wire [39:0]               lrq_user;           // TUSER for request {SrcID,DestID,3'b0,RESPONSE,1'b0,CRF,1'b0}
  wire                      lrq_header_stage;   // Generating the header for a request
  reg                       lrq_data_stage;     // Generating the data for a request
  wire                      lrq_active;         // The lrtx_req interface is active (ready && valid)
  wire                      lrq_sof;            // The lrtx_req interface fisrt beat is accepted by the arb
  wire                      lrq_last;           // The lrtx_req interface last beat is accepted by the arb
  reg                       lrq_last_hold;      // The last active beat was the lastr beat of a packet
  wire                      lrq_rreq_sent;      // A read request was accepted for transmission by the arbiter
  wire                      lrq_wreq_sent;      // A write request was accepted for transmission by the arbiter
  // }}} end Wire Declarations

  // {{{ Register Reset
  // Must register the resets before use to reduce fanout
  always @(posedge log_clk) begin
    log_rst_q   <= #TCQ log_rst;
  end
  // Create an and'ed reset for the maintr logic in order to allow implementation of a link timeout
  // Also re-register the reset - used to set the READY signals
  always @(posedge log_clk) begin
    maintrlog_rst_q   <= #TCQ maintr_rst || log_rst;
    maintrlog_rst_qq  <= #TCQ maintrlog_rst_q;
  end
  // }}} end Register Reset

  // {{{ User Interface - lru
  // + {{{ User Read Interface +
  // Contains the AXI-Lite maint read address channel and read response channel interfaces
  //----------------------------------------
  assign lru_aractive = LR_maintr_arready && UG_maintr_arvalid; // Address is transferred
  assign lru_ractive  = UG_maintr_rready  && LR_maintr_rvalid;  // Response is transferred

  // Register read address on address transfer
  always @(posedge log_clk) begin
    // No reset needed because only sampled when address is valid
    if (lru_aractive) begin
      lru_raddr <= #TCQ UG_maintr_araddr;
    end
  end

  // Create flag indicating that read address has been received
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lru_aractive_q    <= #TCQ 1'b0;
    end else begin
      lru_aractive_q    <= #TCQ lru_aractive;
    end
  end

  // Create the arready signal - should be high until address received, set back high on response xfer
  // Tie low if core can not send MAINT packets and if local config access is unsupported
  always @(posedge log_clk) begin
    if (maintrlog_rst_q) begin
      LR_maintr_arready      <= #TCQ 1'b0;
    end else if (MAINT_SOURCE == 0) begin
      LR_maintr_arready      <= #TCQ 1'b0;
    end else if (maintrlog_rst_qq) begin
      LR_maintr_arready      <= #TCQ 1'b1;
    end else if (lru_ractive) begin
      LR_maintr_arready      <= #TCQ 1'b1;
    end else if (lru_aractive) begin
      LR_maintr_arready      <= #TCQ 1'b0;
    end
  end

  // If there is a read response, register the data and response
  always @(posedge log_clk) begin
    // No reset because these are only valid when LR_maintr_rvalid is asserted
    if (lrm_ur_got_rresp) begin
      LR_maintr_rresp <= #TCQ lrm_ur_rresp;
      LR_maintr_rdata <= #TCQ lrm_ur_rdata;
    end
  end

  // Create the rvalid signal - should be high after response rcvd, cleared on response xfer
  // Tie low if core can not send MAINT packets and if local config access is unsupported
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LR_maintr_rvalid      <= #TCQ 1'b0;
    end else if (MAINT_SOURCE == 0) begin
      LR_maintr_rvalid      <= #TCQ 1'b0;
    end else if (lrm_ur_got_rresp) begin
      LR_maintr_rvalid      <= #TCQ 1'b1;
    end else if (lru_ractive) begin
      LR_maintr_rvalid      <= #TCQ 1'b0;
    end
  end

  //*ASSERTION*
  //(ap_no_lru_aractive_and_ractive): lru_ractive and lru_aractive should not be asserted together
  //(ap_lru_rvalid_set_and_clr): lru_ractive and lrm_ur_got_rresp should not be asserted together
  //(ap_unexpected_lrm_ur_rresp): lrm_ur_got_rresp should not assert if LR_maintr_arready is set

  //IPCV: UG_maintr_rready input used unregistered (to clear rvalid and set arready)
  //IPCV: UG_maintr_arvalid input used unregistered (to clear arready, set got_raddr, and as CE on raddr and ruser)

  // + }}} end User Read Interface +

  // + {{{ User Write Interface +
  // Contains the AXI-Lite maint write address, write data, and write response channel interfaces
  //----------------------------------------
  assign lru_awactive    = LR_maintr_awready && UG_maintr_awvalid; // Address is transferred
  assign lru_wactive     = LR_maintr_wready  && UG_maintr_wvalid;  // Data and Strobe are transferred
  assign lru_bactive     = UG_maintr_bready  && LR_maintr_bvalid;  // Response is transferred

  // Register write address on address transfer
  always @(posedge log_clk) begin
    // No reset because the write address is only sampled on a valid address transfer
    if (lru_awactive) begin
      lru_waddr         <= #TCQ UG_maintr_awaddr;
    end
  end

  // Create flag indicating that write address has been received
  always @(posedge log_clk) begin
    if (maintrlog_rst_q) begin
      lru_got_waddr     <= #TCQ 1'b0;
    end else if (lru_awactive) begin
      lru_got_waddr     <= #TCQ 1'b1;
    end else if (lru_got_waddr && lru_got_wdata) begin
      lru_got_waddr     <= #TCQ 1'b0;
    end
  end

  // Register write data on data transfer
  always @(posedge log_clk) begin
    // No reset because the data and strobe are only sampled on a valid data transfer
    if (lru_wactive) begin
      lru_wdata         <= #TCQ UG_maintr_wdata;
    end
  end

  // Create flag indicating that write data has been received
  always @(posedge log_clk) begin
    if (maintrlog_rst_q) begin
      lru_got_wdata     <= #TCQ 1'b0;
    end else if (lru_wactive) begin
      lru_got_wdata     <= #TCQ 1'b1;
    end else if (lru_got_waddr && lru_got_wdata) begin
      lru_got_wdata     <= #TCQ 1'b0;
    end
  end

  // Create the awready signal - should be high until address received, set back high on response xfer
  // Tie low if core can not send MAINT packets and if local config access is unsupported
  always @(posedge log_clk) begin
    if (maintrlog_rst_q) begin
      LR_maintr_awready  <= #TCQ 1'b0;
    end else if (MAINT_SOURCE == 0) begin
      LR_maintr_awready  <= #TCQ 1'b0;
    end else if (maintrlog_rst_qq) begin
      LR_maintr_awready  <= #TCQ 1'b1;
    end else if (lru_bactive) begin
      LR_maintr_awready  <= #TCQ 1'b1;
    end else if (lru_awactive) begin
      LR_maintr_awready  <= #TCQ 1'b0;
    end
  end

  // Create the wready signal - should be high until data received, set back high on response xfer
  // Tie low if core can not send MAINT packets and if local config access is unsupported
  always @(posedge log_clk) begin
    if (maintrlog_rst_q) begin
      LR_maintr_wready   <= #TCQ 1'b0;
    end else if (MAINT_SOURCE == 0) begin
      LR_maintr_wready   <= #TCQ 1'b0;
    end else if (maintrlog_rst_qq) begin
      LR_maintr_wready   <= #TCQ 1'b1;
    end else if (lru_bactive) begin
      LR_maintr_wready   <= #TCQ 1'b1;
    end else if (lru_wactive) begin
      LR_maintr_wready   <= #TCQ 1'b0;
    end
  end

  // If there is a write response, register it
  always @(posedge log_clk) begin
    // No reset because these are only valid when LR_maintr_bvalid is asserted
    if (lrm_uw_got_wresp) begin
      LR_maintr_bresp    <= #TCQ lrm_uw_wresp;
    end
  end

  // Create the bvalid signal - should be high after response rcvd, cleared on response xfer
  // Tie low if core can not send MAINT packets and if local config access is unsupported
  always @(posedge log_clk) begin
    if (maintrlog_rst_q) begin
      LR_maintr_bvalid   <= #TCQ 1'b0;
    end else if (MAINT_SOURCE == 0) begin
      LR_maintr_bvalid   <= #TCQ 1'b0;
    end else if (lrm_uw_got_wresp) begin
      LR_maintr_bvalid   <= #TCQ 1'b1;
    end else if (lru_bactive) begin
      LR_maintr_bvalid   <= #TCQ 1'b0;
    end
  end

  //*ASSERTION*
  //(ap_no_lru_awactive_and_bactive): lru_bactive and lru_awactive should not be asserted together
  //(ap_no_lru_wactive_and_bactive): lru_bactive and lru_wactive should not be asserted together
  //(ap_lru_bvalid_set_and_clr): lru_bactive and lrm_uw_got_wresp should not be asserted together
  //(ap_unexpected_lrm_uw_wresp): lrm_uw_got_wresp should not assert if LR_maintr_awready or LR_maintr_wready are set

  //*COVERAGE*
  //(cp_got_waddr_and_not_wdata): got_wdata is high and got_waddr is low
  //(cp_got_wdata_and_not_waddr): got_waddr is high and got_wdata is low
  //(cp_awactive_and_wactive): write data and address transferred simultaneously

  //IPCV: UG_maintr_bready input used unregistered (to clear bvalid and set awready and wready)
  //IPCV: UG_maintr_awvalid input used unregistered (to clear awready, set got_waddr, and in CE on waddr and wuser)
  //IPCV: UG_maintr_wvalid input used unregistered (to clear wready, set got_wdata, and in CE on wdata)

  // + }}} end User Write Interface +
  // }}} end User Interface - lru

  // {{{ Arbiter RX Interface - lrr
  // Contains the Arb RX interface and indicates the type of packet being received
  //----------------------------------------
  assign lrr_active  = LR_lrrx_tready && LA_lrrx_tvalid; // Data is transferred

  // Register tlast so that we can find the SOF
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lrr_tlast_hold <=  #TCQ 1'b1; // Reset to one so that sof asserts for the first frame
      lrr_sof_hold   <=  #TCQ 1'b0;
    end else if (lrr_active) begin
      lrr_tlast_hold <=  #TCQ LA_lrrx_tlast;
      lrr_sof_hold   <=  #TCQ lrr_sof;
    end
  end

  // The sof is valid when lrr_tlast_hold is high and there is a data transfer
  assign lrr_sof     = lrr_active && lrr_tlast_hold;

  // Create a flag indicating the last beat of a packet on the lrrx interface
  assign lrr_last    = lrr_active && LA_lrrx_tlast;

  // Pick off header fields (only valid on lrr_tlast_hold && LA_lrrx_tvalid)
  assign lrr_tid     = LA_lrrx_tdata[63:56];
  assign lrr_ftype   = LA_lrrx_tdata[55:52];
  assign lrr_ttype   = LA_lrrx_tdata[51:48];
  assign lrr_prio    = LA_lrrx_tdata[46:45];
  assign lrr_crf     = LA_lrrx_tdata[44];
  assign lrr_size    = LA_lrrx_tdata[43:36];
  assign lrr_ok      =~LA_lrrx_tdata[35];
  // Invert bit 2 of address because of HELLO -> sRIO conversion
  assign lrr_addr    = {LA_lrrx_tdata[23:3], ~LA_lrrx_tdata[2], LA_lrrx_tdata[1:0]};

  // Create registered versions of header fields
  always @(posedge log_clk) begin
    // No reset needed because only sampled on valid data
    if (lrr_sof) begin
      lrr_ok_hold     <=  #TCQ lrr_ok;
      lrr_addr_hold   <=  #TCQ lrr_addr[2];
    end
  end

  // Determine the transaction type on the first frame presented by the arbiter
  // READ REQUEST:
  assign lrr_read  = lrr_tlast_hold && LA_lrrx_tvalid &&
                  (((lrr_ftype == FTYPE_NREAD)  && (LCSBA_SUPPORT == 1)) ||       //NREAD
                   ((lrr_ftype == FTYPE_MAINT)  && (lrr_ttype == TTYPE_MREQR)));  //MREQR

  // WRITE REQUEST:
  assign lrr_write = lrr_tlast_hold && LA_lrrx_tvalid &&
                  (((lrr_ftype == FTYPE_NWRITE) && (LCSBA_SUPPORT == 1)) ||       //NWRITE
                   ((lrr_ftype == FTYPE_NWRITE) && (LCSBA_SUPPORT == 1)) ||       //NWRITE_R
                   ((lrr_ftype == FTYPE_MAINT)  && (lrr_ttype == TTYPE_MREQW)));  //MREQW

  // READ RESPONSE:
  assign lrr_rresp = lrr_tlast_hold && LA_lrrx_tvalid &&
                   ((lrr_ftype == FTYPE_MAINT)  && (lrr_ttype == TTYPE_MRESPR));  //MRESPR

  // WRITE RESPONSE:
  assign lrr_wresp = lrr_tlast_hold && LA_lrrx_tvalid &&
                   ((lrr_ftype == FTYPE_MAINT)  && (lrr_ttype == TTYPE_MRESPW));  //MRESPW

  // Note when a sof specifically belongs to a request packet
  assign lrr_req_sof = lrr_sof && (lrr_read || lrr_write);

  // Create flag indicating request is pending
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lrr_req_pending   <= #TCQ 1'b0;
    end else if (lrr_req_sof) begin
      lrr_req_pending   <= #TCQ 1'b1;
    end else if (lrs_resp_sent || (lrm_ext_no_resp && lrm_ext_cfg_wresp)) begin
      lrr_req_pending   <= #TCQ 1'b0;
    end
  end

  // Set ready when a packet comes in that the log_maint has capacity to process:
  // - For unexpected packet types, just read them off and drop silently
  // - For requests, accept if the user does not have a lock on that transaction type
  // - For responses, accept if the log_maint does not already have the response type available to the user
  assign lrr_set_rdy  = lrr_tlast_hold && LA_lrrx_tvalid && !(lrr_read || lrr_write || lrr_rresp || lrr_wresp) ||
                        (!lrr_req_pending && ((lrr_read  && !lrm_ur_read_lock)  ||
                                              (lrr_write && !lrm_uw_write_lock) ||
                                              (lrr_rresp && !LR_maintr_rvalid && !lrm_ur_got_rresp) ||
                                              (lrr_wresp && !LR_maintr_bvalid && !lrm_uw_got_wresp)));

  // Create tready - only high when a desired packet is on the interface
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LR_lrrx_tready    <= #TCQ 1'b0;
    end else if (lrr_last) begin
      LR_lrrx_tready    <= #TCQ  1'b0;
    end else if (lrr_set_rdy) begin
      LR_lrrx_tready    <= #TCQ  1'b1;
    end
  end

  // INTERNAL COVERAGE AND ASSERTIONS
  //*ASSERTION*
  //(ap_lrr_one_transaction_lrrx): Only one of lrr_read, lrr_write, lrr_rresp, and lrr_wresp can be high
  //(ap_lrr_only_one_req): Should not get a request sof while a request is pending
  //(ap_lrr_only_one_rresp): Should not accept a rresp while an rresp is being presented to the user
  //(ap_lrr_only_one_wresp): Should not accept a wresp while a bresp is being presented to the user
  //(ap_lrr_stall_bt_pkts): Should stall between received packets

  //*COVERAGE*
  //(cp_lrr_ok_d_high_rresp): lrr_ok_d is high for an rresp
  //(cp_lrr_ok_d_high_wresp): lrr_ok_d is high for a wresp
  //(cp_lrr_ok_d_low_rresp): lrr_ok_d is low for an rresp
  //(cp_lrr_ok_d_low_wresp): lrr_ok_d is low for a wresp
  //(cp_req_pending_cleared_by_resp_sent): lrr_req_pending is cleared by a resp being sent
  //(cp_req_pending_cleared_with_no_resp): lrr_req_pending is cleared when a write resp rcvd from CF for NWRITE
  //(cp_read_and_req_pending): lrr_read asserts while req_pending is asserted
  //(cp_write_and_req_pending): lrr_write asserts while req_pending is asserted
  //(cp_rresp_and_maintr_rvalid): lrr_rresp asserts while maintr_rvalid is asserted
  //(cp_wresp_and_maintr_bvalid): lrr_wresp asserts while maintr_bvalid is asserted
  //(cp_lrr_prio_enum): Enumerate lrr_prio on lrr_sof
  //(cp_LR_lrrx_tready_set_and_clr): See the set and clear conditions for tready at the same time.

  // ARB INTERFACE COVERAGE AND ASSERTIONS
  //*ASSERTION*
  //(ap_rx_maint_only_if_no_lcsba_support): Only receive MAINT transactions from arb if LCSBA_SUPPORT == 0
  //(ap_rx_ftypes_2_5_8_only): Only receive transactions with FTYPE 2, 5, and 8 from arb
  //(ap_rx_io_pkts_within_lcsba_8bit_devid): Only receive IO transactions from arb within LCSBA space
  //(ap_rx_io_pkts_within_lcsba_16bit_devid): Only receive IO transactions from arb within LCSBA space
  //(ap_rx_valid_does_not_drop_mid_pkt): Once asserted, LA_lrrx_tvalid stays asserted through tlast

  //*COVERAGE*
  //(cp_rx_all_valid_ftypes): Receive all valid FTYPEs and TTYPEs
  //(cp_lrrx_arb_stalls_mid_packet): arb stalls mid-packet on lrrx
  //(cp_lrrx_arb_stalls_beat1): arb stalls after the first beat on lrrx
  //(cp_lrrx_arb_stalls_beat1_rresp): arb stalls after the first beat on an rresp on lrrx

  // }}} end Arbiter RX Interface - lrr

  // {{{ Configuration Fabric Interface - lrc
  // The Log Maint acts as an AXI-Lite Master to the Config Fabric. It presents
  // reads and writes from the user and the link and waits for the responses.
  //----------------------------------------


  // + {{{ Configuration Fabric Read Interface +

  assign lrc_aractive      = CF_cfgr_arready && LR_cfgr_arvalid; // Address is transferred
  assign lrc_ractive       = LR_cfgr_rready  && CF_cfgr_rvalid;  // Response is transferred

  // Create the LR_cfgr_arvalid signal
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LR_cfgr_arvalid     <= #TCQ 1'b0;
    end else if (lrm_ur_read_cfg || lrm_ext_read_cfg) begin
      LR_cfgr_arvalid     <= #TCQ 1'b1;
    end else if (lrc_aractive) begin
      LR_cfgr_arvalid     <= #TCQ 1'b0;
    end
  end

  // Create the LR_cfgr_araddr signal
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LR_cfgr_araddr      <= #TCQ 24'b0;
    end else if (lrm_ext_read_cfg) begin
      LR_cfgr_araddr      <= #TCQ lrr_addr[23:0];
    end else if (lrm_ur_read_cfg) begin
      LR_cfgr_araddr      <= #TCQ lru_raddr[23:0];
    end
  end

  // Tie ARPROT to 0 since it's unused
  assign LR_cfgr_arprot = 3'b0;

  // Create the LR_cfgr_rready signal
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LR_cfgr_rready      <= #TCQ 1'b0;
    end else if (lrc_aractive) begin
      LR_cfgr_rready      <= #TCQ 1'b1;
    end else if (lrc_ractive) begin
      LR_cfgr_rready      <= #TCQ 1'b0;
    end
  end

  // Register the data and response when the response is transfered
  always @(posedge log_clk) begin
    // No reset needed because only sampled on valid response transfer
    if (lrc_ractive) begin
      lrc_rdata           <= #TCQ CF_cfgr_rdata;
      lrc_rresp           <= #TCQ CF_cfgr_rresp;
    end
  end

  // Indicate when a read response is ready - register to reduce fanout on core input CF_cfgr_rvalid
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lrc_got_rresp       <= #TCQ 1'b0;
    end else begin
      lrc_got_rresp       <= #TCQ lrc_ractive;
    end
  end

  //IPCV: CF_cfgr_rvalid input used unregistered (to register data and resp, to clear rready, and for lrc_got_rresp)
  //IPCV: CF_cfgr_arready input used unregistered (to clear LR_cfgr_arvalid)

  // + }}} end Configuration Fabric Read Interface +

  // + {{{ Configuration Fabric Write Interface +

  assign lrc_awactive      = CF_cfgr_awready && LR_cfgr_awvalid; // Address is transferred
  assign lrc_wactive       = CF_cfgr_wready  && LR_cfgr_wvalid;  // Data is transferred
  assign lrc_bactive       = LR_cfgr_bready  && CF_cfgr_bvalid;  // Response is transferred

  // Create the LR_cfgr_awvalid signal
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LR_cfgr_awvalid     <= #TCQ 1'b0;
    end else if (lrm_uw_write_cfg || lrm_ext_write_cfg) begin
      LR_cfgr_awvalid     <= #TCQ 1'b1;
    end else if (lrc_awactive) begin
      LR_cfgr_awvalid     <= #TCQ 1'b0;
    end
  end

  // Tie AWPROT to 0 since it's unused
  assign LR_cfgr_awprot = 3'b0;

  // Create the LR_cfgr_wvalid signal
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LR_cfgr_wvalid      <= #TCQ 1'b0;
    end else if (lrm_uw_write_cfg || lrm_ext_write_cfg) begin
      LR_cfgr_wvalid      <= #TCQ 1'b1;
    end else if (lrc_wactive) begin
      LR_cfgr_wvalid      <= #TCQ 1'b0;
    end
  end

  // Create the LR_cfgr_wdata signal, using data from arb request or user as appropriate
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LR_cfgr_wdata       <= #TCQ 32'b0;
    end else if (lrm_ext_write_cfg) begin
      LR_cfgr_wdata       <= #TCQ lrr_addr_hold ? LA_lrrx_tdata[31:0] : LA_lrrx_tdata[63:32];
    end else if (lrm_uw_write_cfg) begin
      LR_cfgr_wdata       <= #TCQ lru_wdata;
    end
  end

  // Tie wstrb high because only WORD accesses are allowed - see RapidIO Spec 4.1.10
  assign LR_cfgr_wstrb = 4'hF;

  // Create the LR_cfgr_awaddr signal
  // (on arb request, update awaddr a cycle early to avoid registering it twice)
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LR_cfgr_awaddr      <= #TCQ 24'b0;
    end else if (lrm_ext_got_waddr) begin
      LR_cfgr_awaddr      <= #TCQ lrr_addr;
    end else if (lrm_uw_write_cfg) begin
      LR_cfgr_awaddr      <= #TCQ lru_waddr[23:0];
    end
  end

  // Create the LR_cfgr_bready signal
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LR_cfgr_bready      <= #TCQ 1'b0;
    end else if (lrc_awactive) begin
      LR_cfgr_bready      <= #TCQ 1'b1;
    end else if (lrc_bactive) begin
      LR_cfgr_bready      <= #TCQ 1'b0;
    end
  end

  // Register the response when the response is transfered
  always @(posedge log_clk) begin
    // No reset needed because only sampled on valid response transfer
    if (lrc_bactive) begin
      lrc_wresp           <= #TCQ CF_cfgr_bresp;
    end
  end

  // Signal that a write response is ready
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lrc_got_wresp       <= #TCQ 1'b0;
    end else begin
      lrc_got_wresp       <= #TCQ lrc_bactive;
    end
  end


  // CONFIG FABRIC INTERFACE COVERAGE AND ASSERTIONS
  //*COVERAGE*
  //(cp_cfgr_waddr_before_wdata): The waddr is accepted before the wdata
  //(cp_cfgr_wdata_before_waddr): The wdata is accepted before the waddr

  //IPCV: CF_cfgr_bvalid input used unregistered (to register resp, to clear bready, and for lrc_got_wresp)
  //IPCV: CF_cfgr_awready input used unregistered (to clear LR_cfgr_awvalid)
  //IPCV: CF_cfgr_wready input used unregistered (to clear LR_cfgr_wvalid)

  // + }}} end Configuration Fabric Write Interface +
  // }}} end Configuration Fabric Interface - lrc

  // {{{ Maint Request Info Register - lri
  // This configuration register stored in the LOG Maint allows users to set
  // the Destination ID, TID, prio, CRF, and VC fields for outgoing maintenance
  // requests.
  //----------------------------------------

  // Capture writes to Request Info Register (except TID field which is handled below)
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lri_req_vc              <= #TCQ 1'b0;
      lri_req_prio            <= #TCQ 2'b01;
      lri_req_crf             <= #TCQ 1'b0;
      lri_req_destid          <= #TCQ 16'b0;
    // Update on user write
    end else if (lrm_uw_info_reg_wen) begin
      lri_req_vc            <= #TCQ (VC == 1) ? lru_wdata[19] : 1'b0;
      lri_req_prio          <= #TCQ lru_wdata[18:17];
      lri_req_crf           <= #TCQ (CRF_SUPPORT == 1) ? lru_wdata[16] : 1'b0;
      lri_req_destid[15:8]  <= #TCQ lru_wdata[15:8];
      lri_req_destid[7:0]   <= #TCQ lru_wdata[7:0];
    // Update on external write
    end else if (lrm_ext_info_reg_wen) begin
      lri_req_vc            <= #TCQ (VC == 1) ? LA_lrrx_tdata[51] : 1'b0;
      lri_req_prio          <= #TCQ LA_lrrx_tdata[50:49];
      lri_req_crf           <= #TCQ (CRF_SUPPORT == 1) ? LA_lrrx_tdata[48] : 1'b0;
      lri_req_destid[15:8]  <= #TCQ LA_lrrx_tdata[47:40];
      lri_req_destid[7:0]   <= #TCQ LA_lrrx_tdata[39:32];
    end
  end

  // Compute the next tid to be used for an outgoing MREQ
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lri_req_next_tid  <= #TCQ 8'b0;
    end else if (lrm_uw_info_reg_wen) begin
      lri_req_next_tid  <= #TCQ lru_wdata[31:24];
    // Load the written value on a write
    end else if (lrm_ext_info_reg_wen) begin
      lri_req_next_tid  <= #TCQ LA_lrrx_tdata[63:56];
    // Increment when a new request is formed
    end else if (lrq_start) begin
      lri_req_next_tid  <= #TCQ lri_req_next_tid + 1'b1;
    end
  end

                                                        // core  (spec)   Description
                                                        // ----------------------------
  // Maintenance Request Information CSR
  assign lri_csr_lr_000  = {lri_req_next_tid,           // 31:24  (0:7)   TID for next outgoing MREQ
                            4'b0,                       // 23:20  (8:11)  Reserved
                            lri_req_vc,                 // 19     (12)    VC for outgoing MREQs
                            lri_req_prio,               // 18:17  (13:14) Prio for outgoing MREQs
                            lri_req_crf,                // 16     (15)    CRF for outgoing MREQs
                            lri_req_destid};            // 15:0   (16:31) Destination Device ID for outgoing MREQs

  //*COVERAGE*
  //(cp_lri_req_next_tid_rolls_over): The next TID counter rolls over
  //(cp_lri_req_next_tid_load_local): The next TID counter is loaded with a new TID from a local write
  //(cp_lri_req_next_tid_load_ext): The next TID counter is loaded with a new TID from an external write
  //(cp_lrm_uw_info_reg_wen): The Maint Request Info Register is written by the user
  //(cp_lrm_ext_info_reg_wen): The Maint Request Info Register is written by the remote device
  //(cp_tid_increments_sending_request): The Maint Request Info Register is incremented when a request is sent

  //*CROSS*
  //(cr_tid_updates): each combination of tid update mechanisms occurs

  // }}} end Maint Request Info Register - lri

  // {{{ Read and Write Managers - lrm
  // The read and write managers are responsible for tracking the phase of
  // each transaction and creating flags to other blocks when action is needed.
  //----------------------------------------

  // + {{{ User Read Manager - lrm_ur +
  // The User Read Manager is responsible for completing user reads. For local
  // reads, it waits until the config fabric is ready then forwards the read
  // there. For remote reads, it signals the packet generator to form a read
  // for transmit on the link, then monitors incoming read responses and
  // returns the response to the user when the TID matches the read request.
  // It also implements a port timeout counter for remote reads.
  //----------------------------------------

  // Create a signal indicating the type of read when one is available
  assign lrm_ur_info      = (!(|lru_raddr[31:24]) && (lru_raddr[23:2] == CSR_INFO_REG[23:2]));
  assign lrm_ur_local     = (!(|lru_raddr[31:24]) && !lrm_ur_info);
  assign lrm_ur_remote    =   (|lru_raddr[31:24]);

  // Create a signal indicating that a read is pending
  always @(posedge log_clk) begin
    if (maintrlog_rst_q) begin
      lrm_ur_info_pend    <= #TCQ 1'b0;
      lrm_ur_local_pend   <= #TCQ 1'b0;
      lrm_ur_remote_pend  <= #TCQ 1'b0;
    end else if (lrm_ur_got_rresp) begin
      lrm_ur_info_pend    <= #TCQ 1'b0;
      lrm_ur_local_pend   <= #TCQ 1'b0;
      lrm_ur_remote_pend  <= #TCQ 1'b0;
    end else if (lru_aractive_q) begin
      lrm_ur_info_pend    <= #TCQ lrm_ur_info;
      lrm_ur_local_pend   <= #TCQ lrm_ur_local;
      lrm_ur_remote_pend  <= #TCQ lrm_ur_remote;
    end
  end

  // Create a lock signal to indicate when the User Read Manager "owns" the CF read channels
  always @(posedge log_clk) begin
    if (maintrlog_rst_q) begin
      lrm_ur_read_lock    <= #TCQ 1'b0;
    end else if (LR_maintr_rvalid) begin
      lrm_ur_read_lock    <= #TCQ 1'b0;
    // Link reads have higher priority, so check that none are queued up
    end else if (lrm_ur_local_pend && !lrr_read && !lrm_ext_read_lock) begin
      lrm_ur_read_lock    <= #TCQ 1'b1;
    end
  end

  // Create a registered version of the lock signal so that the rising edge can be detected
  always @(posedge log_clk) begin
    if (maintrlog_rst_q) begin
      lrm_ur_read_lock_q  <= #TCQ 1'b0;
    end else begin
      lrm_ur_read_lock_q  <= #TCQ lrm_ur_read_lock;
    end
  end

  // Create a signal to use to set LR_cfgr_arvalid when a user read has arrived and the user "owns" the interface
  assign lrm_ur_read_cfg = lrm_ur_read_lock && !lrm_ur_read_lock_q;

  // Signal to the Packet Generator to create a read request
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lrm_ur_rreq_gen    <= #TCQ 1'b0;
    end else if (lru_aractive_q && lrm_ur_remote) begin
      lrm_ur_rreq_gen    <= #TCQ 1'b1;
    end else if (lrq_rreq_sent) begin
      lrm_ur_rreq_gen    <= #TCQ 1'b0;
    end
  end

  // Create hopcount for use in request generator
  assign lrm_ur_hopcount = lru_raddr[31:24] - 1'b1;

  // Save the TID used on the outgoing request
  always @(posedge log_clk) begin
    if (maintrlog_rst_q) begin
      lrm_ur_tid      <= #TCQ 8'b0;
    end else if (lrq_start && (lrq_pktsel == SENDING_READ)) begin
      lrm_ur_tid      <= #TCQ lri_req_next_tid;
    end
  end

  // Check TID of incoming response (only used after rresp is received from link partner)
  always @(posedge log_clk) begin
    if (maintrlog_rst_q) begin
      lrm_ur_tid_match   <= #TCQ 1'b0;
    end else if (lrr_last) begin
      lrm_ur_tid_match   <= #TCQ 1'b0;
    end else if (lrm_ur_remote_pend && lrr_rresp && lrr_sof && (lrr_tid == lrm_ur_tid)) begin
      lrm_ur_tid_match   <= #TCQ 1'b1;
    end
  end

  // Create flag when response is available
  assign lrm_ur_got_rresp = (lrm_ur_remote_pend && lrm_ur_tid_match && lrr_last)  || // TID match on response
                             lrm_ur_info_pend                                     || // Read to Request Info register
                            (lrm_ur_read_lock && lrc_got_rresp);                     // Response rcvd from local CFG

  // Create Response
  assign lrm_ur_rresp     = lrm_ur_remote_pend ? {!lrr_ok_hold, 1'b0} :
                            lrm_ur_info_pend   ? 2'b0                                     :
                                            lrc_rresp;
  // Create read data
  assign lrm_ur_rdata     = lrm_ur_remote_pend ? (lru_raddr[2] ? LA_lrrx_tdata[31:0] : LA_lrrx_tdata[63:32]) :
                            lrm_ur_info_pend   ?  lri_csr_lr_000                                             :
                                             lrc_rdata;

  //*COVERAGE*
  //(cp_local_rresp_rcvd): A response is received from the CF for a local read

  // + }}} end User Read Manager - lrm_ur +

  // + {{{ User Write Manager - lrm_uw +
  // The User Write Manager is responsible for completing user writes. For
  // local writes, it waits until the config fabric is ready then forwards the
  // write there. For remote writes, it signals the packet generator to form a
  // write for transmit on the link, then monitors incoming write responses and
  // returns the response to the user when the TID matches the write request.
  // It also implements a port timeout counter for remote writes.
  //----------------------------------------


  // Create a signal indicating the type of write when one is available
  assign lrm_uw_info    = !(|lru_waddr[31:24]) && (lru_waddr[23:2] == CSR_INFO_REG[23:2]);
  assign lrm_uw_local   = !(|lru_waddr[31:24]) && !lrm_uw_info;
  assign lrm_uw_remote  =  (|lru_waddr[31:24]);

  // Create a signal indicating that the type of write that is pending
  always @(posedge log_clk) begin
    if (maintrlog_rst_q) begin
      lrm_uw_info_pend      <= #TCQ 1'b0;
      lrm_uw_local_pend     <= #TCQ 1'b0;
      lrm_uw_remote_pend    <= #TCQ 1'b0;
    end else if (lrm_uw_got_wresp) begin
      lrm_uw_info_pend      <= #TCQ 1'b0;
      lrm_uw_local_pend     <= #TCQ 1'b0;
      lrm_uw_remote_pend    <= #TCQ 1'b0;
    end else if (lru_got_waddr && lru_got_wdata) begin
      lrm_uw_info_pend      <= #TCQ lrm_uw_info;
      lrm_uw_local_pend     <= #TCQ lrm_uw_local;
      lrm_uw_remote_pend    <= #TCQ lrm_uw_remote;
    end
  end

  // Create a lock signal to indicate when the User Write Manager "owns" the CF write channels
  always @(posedge log_clk) begin
    if (maintrlog_rst_q) begin
      lrm_uw_write_lock     <= #TCQ 1'b0;
    end else if (LR_maintr_bvalid) begin
      lrm_uw_write_lock     <= #TCQ 1'b0;
    // Link writes have higher priority, so check that none are queued up and there are none in progress
    end else if (lrm_uw_local_pend && !lrr_write && !lrm_ext_write_lock) begin
      lrm_uw_write_lock     <= #TCQ 1'b1;
    end
  end

  // Create a registered version of the lock signal so that the rising edge can be detected
  always @(posedge log_clk) begin
    if (maintrlog_rst_q) begin
      lrm_uw_write_lock_q   <= #TCQ 1'b0;
    end else begin
      lrm_uw_write_lock_q   <= #TCQ lrm_uw_write_lock;
    end
  end

  // Create a signal to use to set LR_cfgr_arvalid when a user write has arrived and the user "owns" the interface
  assign lrm_uw_write_cfg  = lrm_uw_write_lock && !lrm_uw_write_lock_q;

   // Write to the Maintenance Request Info Register
  always @(posedge log_clk) begin
    if (maintrlog_rst_q) begin
      lrm_uw_info_reg_wen   <= #TCQ 1'b0;
    end else begin
      lrm_uw_info_reg_wen   <= #TCQ lru_got_wdata && lru_got_waddr && lrm_uw_info;
    end
  end

  // Signal to the Packet Generator to create a write request
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lrm_uw_wreq_gen       <= #TCQ 1'b0;
    end else if (lru_got_wdata && lru_got_waddr && lrm_uw_remote) begin
      lrm_uw_wreq_gen       <= #TCQ 1'b1;
    end else if (lrq_wreq_sent) begin
      lrm_uw_wreq_gen       <= #TCQ 1'b0;
    end
  end

  // Save the TID used on the outgoing request
  always @(posedge log_clk) begin
    if (maintrlog_rst_q) begin
      lrm_uw_tid      <= #TCQ 8'b0;
    end else if (lrq_start && (lrq_pktsel == SENDING_WRITE)) begin
      lrm_uw_tid      <= #TCQ lri_req_next_tid;
    end
  end

  // Create hopcount for use in request generator
  assign lrm_uw_hopcount = lru_waddr[31:24] - 1'b1;

  // Check TID of incoming response
  always @(posedge log_clk) begin
    if (maintrlog_rst_q) begin
      lrm_uw_tid_match <= #TCQ 1'b0;
    end else begin
      lrm_uw_tid_match <= #TCQ lrm_uw_remote_pend && lrr_wresp && lrr_sof && (lrr_tid == lrm_uw_tid);
    end
  end

  // Create flag when response is available
  assign lrm_uw_got_wresp  = (lrm_uw_remote_pend && lrm_uw_tid_match) ||  // Response rcvd from link partner
                              lrm_uw_info_reg_wen                     ||  // Write to Req Info reg (assume complete)
                             (lrm_uw_write_lock && lrc_got_wresp);        // Response rcvd from local CFG

  // Create Response
  assign lrm_uw_wresp      = lrm_uw_local_pend ? lrc_wresp :
                             lrm_uw_info_pend  ? 2'b0      :
                             {!lrr_ok_hold, 1'b0};

  //*COVERAGE*
  //(cp_early_wresp_bad_strobe): An early response is returned for a remote write due to an invalid strobe
  //(cp_local_wresp_rcvd): A response is received from the CF for a local write

  // + }}} end User Write Manager - lrm_uw +

  // + {{{ External Request Manager - lrm_ext +
  // The External Request Manager is responsible for completing requests from
  // the link partner. It checks the size and waits until the config fabric is
  // ready, then forwards the request there. When the response is available, it
  // signals the response generator to form the appropriate response for transmit
  // on the link (if a response is required based on the request type).
  //----------------------------------------

  // The lrm_ext_read_lock signal indicates that the link read manager "owns" the CF read interface
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lrm_ext_read_lock   <= #TCQ 1'b0;
    end else if (lrs_resp_sent) begin
      lrm_ext_read_lock   <= #TCQ 1'b0;
    end else if (lrr_read && !lrm_ur_read_lock && !lrr_req_pending) begin
      lrm_ext_read_lock   <= #TCQ 1'b1;
    end
  end

  // The lrm_ext_write_lock signal indicates that the external write manager "owns" the CF write interface
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lrm_ext_write_lock  <= #TCQ 1'b0;
    end else if (lrs_resp_sent || (lrm_ext_no_resp && lrm_ext_cfg_wresp)) begin
      lrm_ext_write_lock  <= #TCQ 1'b0;
    end else if (lrr_write && !lrm_uw_write_lock && !lrr_req_pending) begin
      lrm_ext_write_lock  <= #TCQ 1'b1;
    end
  end

  // A read/write is ready if an external read/write is in progress (locked) and the last signal is asserted by the arb
  assign lrm_ext_read_rdy  = lrr_last && lrm_ext_read_lock;
  assign lrm_ext_write_rdy = lrr_last && lrm_ext_write_lock;

  // Check that the read is no larger than 4 bytes and has a valid TTYPE
  assign lrm_ext_size_ok    = (lrr_size < 8'h04);
  assign lrm_ext_type_ok    = (((lrr_ftype == FTYPE_NWRITE) && (lrr_ttype == TTYPE_NWRITE))   ||
                               ((lrr_ftype == FTYPE_NWRITE) && (lrr_ttype == TTYPE_NWRITE_R)) ||
                               ((lrr_ftype == FTYPE_NREAD)  && (lrr_ttype == TTYPE_NREAD))    ||
                               // Do not need to check ttype on MAINT b/c already checked in lrr_read/lrr_write
                                (lrr_ftype == FTYPE_MAINT));
  assign lrm_ext_req_ok     = lrm_ext_size_ok && lrm_ext_type_ok;

  // Check whether the request has valid size/TTYPE, whether it requires a response, and whether it's I/O or MAINT
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lrm_ext_req_ok_hold <= #TCQ 1'b0;
      lrm_ext_no_resp     <= #TCQ 1'b0;
    end else if (lrr_req_sof) begin
      lrm_ext_req_ok_hold <= #TCQ lrm_ext_req_ok;
      lrm_ext_no_resp     <= #TCQ (LCSBA_SUPPORT == 1) && (lrr_ftype == FTYPE_NWRITE) && (lrr_ttype == TTYPE_NWRITE);
    end
  end

  // Once a read is ready, present it to the Cfg Fabric Interface or request an error response
  assign lrm_ext_info_reg_ren  = lrm_ext_read_rdy &&  lrm_ext_req_ok && (lrr_addr[23:2] == CSR_INFO_REG[23:2]);
  assign lrm_ext_read_cfg      = lrm_ext_read_rdy &&  lrm_ext_req_ok && !lrm_ext_info_reg_ren;
  assign lrm_ext_read_err      = lrm_ext_read_rdy && !lrm_ext_req_ok;

  // If the read is to the Request Info register, set a flag so that the proper read data is used in the response
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lrm_ext_info_read     <= #TCQ 1'b0;
    end else if (lrs_resp_sent) begin
      lrm_ext_info_read     <= #TCQ 1'b0;
    end else if (lrm_ext_info_reg_ren) begin
      lrm_ext_info_read     <= #TCQ 1'b1;
    end
  end

  // To avoid registering the write address an extra time, create a flag used to overwrite the addr to the CF on beat 2
  assign lrm_ext_got_waddr  = lrm_ext_write_lock && lrr_sof;

  // When an incoming write is targeted to the Maintenance Request Info register, create a write enable
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lrm_ext_info_reg_write  <= #TCQ 1'b0;
    end else if ((lrr_addr[23:2] == CSR_INFO_REG[23:2]) && lrm_ext_got_waddr) begin
      lrm_ext_info_reg_write  <= #TCQ 1'b1;
    end else if (lrm_ext_write_rdy) begin
      lrm_ext_info_reg_write  <= #TCQ 1'b0;
    end
  end

  // Once a write is ready, present it to the Cfg Fabric Interface or request an error response
  assign lrm_ext_info_reg_wen = lrm_ext_write_rdy &&  lrm_ext_info_reg_write &&  lrm_ext_req_ok_hold;
  assign lrm_ext_write_cfg    = lrm_ext_write_rdy && !lrm_ext_info_reg_wen   &&  lrm_ext_req_ok_hold;
  assign lrm_ext_write_err    = lrm_ext_write_rdy && !lrm_ext_info_reg_wen   && !lrm_ext_req_ok_hold;


  // A response on the Cfg Fabric interface is ours if the lock signal is asserted
  assign lrm_ext_cfg_rresp  = lrc_got_rresp && lrm_ext_read_lock;
  assign lrm_ext_cfg_wresp  = lrc_got_wresp && lrm_ext_write_lock;

  // Select the response FTYPE and TTYPE - only valid on lrr_req_sof
  always @* begin
    case(lrr_ftype)
      FTYPE_NWRITE: begin
        lrm_ext_resp_ftype  = (lrr_ttype == TTYPE_NWRITE) ? 4'bx : FTYPE_RESP;
        lrm_ext_resp_ttype  = (lrr_ttype == TTYPE_NWRITE) ? 4'bx : TTYPE_RESPW;
      end
      FTYPE_NREAD: begin
        lrm_ext_resp_ftype  = FTYPE_RESP;
        lrm_ext_resp_ttype  = TTYPE_RESPR;
      end
      FTYPE_MAINT: begin
        lrm_ext_resp_ftype  = FTYPE_MAINT;
        lrm_ext_resp_ttype  = (lrr_ttype == TTYPE_MREQR) ? TTYPE_MRESPR : TTYPE_MRESPW;
      end
      default:     begin
        lrm_ext_resp_ftype  = 4'bx;
        lrm_ext_resp_ttype  = 4'bx;
      end
    endcase
  end

  // Increment priority for response - only valid on lrr_req_sof
  assign lrm_ext_resp_prio = lrr_prio == 2'b11 ? 2'b11 : lrr_prio + 2'b01;

  // Create the response status (4'b0000 - OK/done, 4'b0111 - Error)
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lrm_ext_resp_err  <= #TCQ 1'b0;
    end else if (lrm_ext_info_reg_wen || lrm_ext_info_reg_ren) begin //Assume pass if targeting Req Info reg
      lrm_ext_resp_err  <= #TCQ 1'b0;
    end else if (lrm_ext_cfg_wresp) begin
      lrm_ext_resp_err  <= #TCQ |lrc_wresp;
    end else if (lrm_ext_cfg_rresp) begin
      lrm_ext_resp_err  <= #TCQ |lrc_rresp;
    end else if (lrm_ext_read_err || lrm_ext_write_err) begin
      lrm_ext_resp_err  <= #TCQ 1'b1;
    end
  end

  // Request a response for a bad read or when a response is received from the Cfg Fabric
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lrm_ext_rresp_gen   <= #TCQ 1'b0;
    end else if (lrs_resp_sent) begin
      lrm_ext_rresp_gen   <= #TCQ 1'b0;
    end else if (lrm_ext_read_err || lrm_ext_cfg_rresp || lrm_ext_info_reg_ren) begin
      lrm_ext_rresp_gen   <= #TCQ 1'b1;
    end
  end

  // Request a response for a bad write, when a response is received from the Cfg Fabric, or after a Req Info write
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lrm_ext_wresp_gen   <= #TCQ 1'b0;
    end else if (lrs_resp_sent || (lrm_ext_no_resp && lrm_ext_cfg_wresp)) begin
      lrm_ext_wresp_gen   <= #TCQ 1'b0;
    end else if (lrm_ext_write_err || lrm_ext_cfg_wresp || lrm_ext_info_reg_wen) begin
      lrm_ext_wresp_gen   <= #TCQ 1'b1;
    end
  end


  //*ASSERTION*
  //(ap_resp_stat_enables_onehot0): The enables for lrm_ext_resp_err are exclusive
  //(ap_write_locks_exclusive): lrm_uw_write_lock and lrm_ext_write_lock should not be high at the same time
  //(ap_read_locks_exclusive): lrm_ur_read_lock and lrm_ext_read_lock should not be high at the same time
  //(ap_ext_locks_exclusive): lrm_ext_write_lock and lrm_ext_read_lock should not be high at the same time
  //(ap_no_resp_req_for_nwrite): lrm_ext_wresp_gen does not assert if lrm_ext_no_resp is high

  //*COVERAGE*
  //(cp_resp_sent_and_lrr_write): lrs_resp_sent and lrr_write are both high
  //(cp_resp_sent_and_lrr_read): lrs_resp_sent and lrr_read are both high
  //(cp_lrm_ext_resp_prio_enum): enumerate lrm_ext_resp_prio on lrr_sof
  //(cp_lrm_ext_read_err_high): lrm_ext_read_err is high
  //(cp_lrm_ext_write_err_high): lrm_ext_write_err is high
  //(cp_lrm_ext_info_reg_ren_high): lrm_ext_info_reg_ren is high
  //(cp_lrm_ext_info_reg_wen_high): lrm_ext_info_reg_wen is high
  //(cp_lrr_read_and_lrm_ur_read_lock): lrr_read and lrm_ur_read_lock are high
  //(cp_lrr_write_and_lrm_uw_write_lock): lrr_write and lrm_uw_write_lock are high
  //(cp_lrm_ext_no_resp_and_lrm_ext_cfg_wresp): wresp rcvd from CF while lrm_ext_no_resp is high
  //(cp_lrm_ext_read_size_err): Read with invalid size detected
  //(cp_lrm_ext_read_type_err): Read with invalid type detected
  //(cp_lrm_ext_write_size_err): Write with invalid size detected
  //(cp_lrm_ext_write_type_err): Write with invalid type detected

  // + }}} end External Request Manager - lrm_ext +
  // }}} end Read and Write Managers - lrm

  // {{{ Arbiter Response Interface - lrs
  // Create responses to send to link partner
  //----------------------------------------

  // The response information is valid if there's a response request and the response wasn't just sent
  assign lrs_valid = (lrm_ext_rresp_gen && !lrs_resp_sent) || (lrm_ext_wresp_gen && !lrs_resp_sent);

  // Determine whether response will have data (only for unerrored reads)
  assign lrs_resp_w_data  = lrm_ext_rresp_gen && !lrm_ext_resp_err;

  // Keep track of which information the Arb TX interface needs
  assign lrs_header_stage = lrs_valid && !lrs_data_stage;

  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lrs_data_stage  <= #TCQ 1'b0;
    end else if (lrs_header_stage && lrs_resp_w_data && lrs_active) begin
      lrs_data_stage  <= #TCQ 1'b1;
    end else if (lrs_data_stage && lrs_active) begin
      lrs_data_stage  <= #TCQ 1'b0;
    end
  end

  assign lrs_active       = LR_lrtx_resp_tvalid && LA_lrtx_resp_tready; // Information is transferred on lrtx_resp

  // Indicate when response has finished sending
  assign lrs_resp_sent    = lrs_active && LR_lrtx_resp_tlast;

  // Form the TDATA output
  always @(posedge log_clk) begin
    if (lrs_header_stage && lrs_active) begin
      // Capture the data on the data stage of a response
      LR_lrtx_resp_tdata          <= #TCQ lrm_ext_info_read ? {lri_csr_lr_000, 32'b0} : {2{lrc_rdata}};
    end else begin
      // Capture the header fields on sof of the request so that they don't have to be double-registered
      if (lrr_req_sof) begin
        LR_lrtx_resp_tdata[63:36] <= #TCQ {lrr_tid,lrm_ext_resp_ftype,lrm_ext_resp_ttype,
                                           1'b0,lrm_ext_resp_prio,lrr_crf,8'b0};
        LR_lrtx_resp_tdata[34:0]  <= #TCQ {1'b0,2'b0,8'hFF,24'b0};
      end
      // Capture the error bit when the response is ready
      if (lrs_header_stage) begin
        LR_lrtx_resp_tdata[35]    <= #TCQ lrm_ext_resp_err;
      end
    end
  end

  // Create the user field based on received values
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LR_lrtx_resp_tuser  <= #TCQ 40'b0;
    end else if (lrr_req_sof) begin
      LR_lrtx_resp_tuser  <= #TCQ {LA_lrrx_tuser[23:8], LA_lrrx_tuser[39:24], 2'b0, 1'b1, 1'b1, 1'b0, LA_lrrx_tuser[2:1], 1'b0};
    end
  end

  // Form the TLAST output
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LR_lrtx_resp_tlast   <= #TCQ 1'b0;
    end else begin
      LR_lrtx_resp_tlast   <= #TCQ !lrs_resp_w_data || lrs_data_stage || (lrs_header_stage && lrs_active);
    end
  end

  // The TKEEP output is always 8'hFF because the interface necessarily uses HELLO format
  assign LR_lrtx_resp_tkeep   = 8'hFF;

  // Register the valid signal to create the valid output
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LR_lrtx_resp_tvalid   <= #TCQ 1'b0;
    end else begin
      LR_lrtx_resp_tvalid   <= #TCQ lrs_valid;
    end
  end

  // INTERNAL COVERAGE AND ASSERTIONS
  //*ASSERTION*
  //(ap_header_data_stage_onehot0): lrs_header_stage, lrs_data_stage, and lrr_req_sof are onehot0

  // ARB INTERFACE COVERAGE AND ASSERTIONS
  //*ASSERTION*
  //(ap_tx_write_resp_1_dword): LOG MAINT only transmits write responses of 1 DWORD
  //(ap_tx_read_resp_1_or_2_dwords): LOG MAINT does not transmit >2 DWORD read response
  //(ap_tx_2_dword_read_resp_ok_status): Read responses of 2 DWORDS have OK status
  //(ap_tx_1_dword_read_resp_err_status): Read responses of 1 DWORDS have ERR status
  //(ap_tx_resp_valid_does_not_drop_mid_pkt): LOG Maint does not deassert tvalid mid-packet
  //(ap_tx_resp_no_b2b): LOG Maint does not issue back-to-back responses

  //*COVERAGE*
  //(cp_tx_err_maint_read_resp): LOG_MAINT transmits a MAINT read response with error status
  //(cp_tx_ok_maint_read_resp): LOG_MAINT transmits a MAINT read response with done status
  //(cp_tx_err_maint_write_resp): LOG_MAINT transmits a MAINT write response with error status
  //(cp_tx_ok_maint_write_resp): LOG_MAINT transmits a MAINT write response with done status
  //(cp_tx_err_io_read_resp): LOG_MAINT transmits an IO read response with error status
  //(cp_tx_ok_io_read_resp): LOG_MAINT transmits an IO read response with done status
  //(cp_tx_err_io_write_resp): LOG_MAINT transmits an IO write response with error status
  //(cp_tx_ok_io_write_resp): LOG_MAINT transmits an IO write response with done status
  //(cp_tx_resp_stalls_mid_packet): arb stalls mid-packet on response
  //(cp_tx_resp_stalls_beat1): arb stalls first beat on response

  // }}} end Arbiter Response Interface - lrs

  // {{{ Arbiter Request Interface - lrq
  // Create requests to send to link partner
  //----------------------------------------

  assign lrq_valid  = (lrm_ur_rreq_gen && !lrq_rreq_sent) || (lrm_uw_wreq_gen && !lrq_wreq_sent);
  assign lrq_start  = lrq_valid && !LR_lrtx_req_tvalid;

  // Select the next packet type. Reads have highest priority.
  assign lrq_pktsel =  (lrm_ur_rreq_gen && !lrq_rreq_sent) ? SENDING_READ  :
                       (lrm_uw_wreq_gen && !lrq_wreq_sent) ? SENDING_WRITE :
                                                             SENDING_NONE  ;

  // Hold the pktsel value so that we know throughout the packet which type was selected
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lrq_pktsel_hold  <= #TCQ SENDING_NONE;
    end else if (lrq_start) begin
      lrq_pktsel_hold  <= #TCQ lrq_pktsel;
    end
  end

  // Select the TTYPE, size, and hopcount for the request based on which packet type is selected
  assign lrq_ttype    = (lrq_pktsel == SENDING_READ) ? TTYPE_MREQR : TTYPE_MREQW;
  assign lrq_size     = 8'h03;
  assign lrq_hopcount = (lrq_pktsel == SENDING_READ) ? lrm_ur_hopcount : lrm_uw_hopcount;
  assign lrq_addr     = (lrq_pktsel == SENDING_READ) ? {lru_raddr[23:3],~lru_raddr[2],2'b0} :
                                                       {lru_waddr[23:3],~lru_waddr[2],2'b0} ;

  // Form packet header
  //FIXVC - Add VC bit when support is added
  assign lrq_header   = {lri_req_next_tid, FTYPE_MAINT, lrq_ttype, 1'b0, lri_req_prio, lri_req_crf,
                         lrq_size, 4'b0, lrq_hopcount, lrq_addr};

  // Form packet data (only used for writes)
  assign lrq_data     = {2{lru_wdata}};

  // Create user signal
  assign lrq_user     = {LC_deviceid, lri_req_destid, 8'h20};

  // Create the data and tlast signals based on the header/data_stage signals
  always @(posedge log_clk) begin
    // No reset needed because only sampled when valid
    if (lrq_active && !LR_lrtx_req_tlast) begin
      LR_lrtx_req_tdata   <= #TCQ lrq_data;
      LR_lrtx_req_tlast   <= #TCQ 1'b1;
    end else if (lrq_start) begin
      LR_lrtx_req_tdata   <= #TCQ lrq_header;
      LR_lrtx_req_tlast   <= #TCQ (lrq_pktsel == SENDING_READ) ? 1'b1 : 1'b0;
    end
  end

  // Register TUSER for arbiter on first valid beat
  always @(posedge log_clk) begin
    // No reset needed because only sampled when valid
    if (lrq_start) begin
      LR_lrtx_req_tuser   <= #TCQ lrq_user;
    end
  end

  assign LR_lrtx_req_tkeep = 8'hFF; // TKEEP is always 8'hFF for HELLO format

  // Create  request valid signal for arbiter
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      LR_lrtx_req_tvalid   <= #TCQ 1'b0;
    end else if (MAINT_SOURCE == 0) begin
      LR_lrtx_req_tvalid   <= #TCQ 1'b0;
    end else begin
      // Enforce a pause between packets so that TID increments appropriately
      LR_lrtx_req_tvalid   <= #TCQ lrq_valid && !(LR_lrtx_req_tlast && lrq_active);
    end
  end

  // Hold the last signal so that the sof can be detected for incrementing the TID
  always @(posedge log_clk) begin
    if (log_rst_q) begin
      lrq_last_hold  <= #TCQ 1'b1; //Reset to 1 so sof is asserted on first packet
    end else if (lrq_active) begin
      lrq_last_hold  <= #TCQ LR_lrtx_req_tlast;
    end
  end

  assign lrq_active        = LR_lrtx_req_tvalid && LA_lrtx_req_tready; // Information is transferred to arb
  assign lrq_sof           = lrq_active && lrq_last_hold;              // First beat of packet is transferred to arb
  assign lrq_last          = lrq_active && LR_lrtx_req_tlast;          // Last beat of packet is transferred to arb

  // Indicate to User Manager that request has been sent
  assign lrq_rreq_sent     = lrq_last && (lrq_pktsel_hold == SENDING_READ);
  assign lrq_wreq_sent     = lrq_last && (lrq_pktsel_hold == SENDING_WRITE);

  // INTERNAL COVERAGE AND ASSERTIONS
  //*COVERAGE*
  //(cp_wreq_and_rreq_gen_rise): lrm_uw_wreq_gen and lrm_ur_rreq_gen rise at the same time
  //(cp_wreq_gen_after_rreq_gen): lrm_uw_wreq_gen rises while lrm_ur_rreq_gen is high
  //(cp_rreq_gen_after_wreq_gen): lrm_ur_rreq_gen rises while lrm_uw_wreq_gen is high
  //(cp_wreq_gen_with_rreq_sent): lrm_uw_wreq_gen rises with lrq_rreq_sent
  //(cp_rreq_gen_with_wreq_sent): lrm_ur_rreq_gen rises with lrq_wreq_sent

  // ARB INTERFACE COVERAGE AND ASSERTIONS
  //*ASSERTION*
  //(ap_tx_mreqw_2_dwords): LOG MAINT only transmits write MREQs of 2 DWORDs
  //(ap_tx_mreqr_1_dwords): LOG MAINT only transmits read MREQs of 1 DWORD
  //(ap_tx_req_valid_does_not_drop_mid_pkt): LOG Maint does not deassert tvalid mid-packet
  //(ap_tx_no_req_if_unsupported): LOG MAINT does not transmit a request if MAINT_SOURCE = 0
  //(ap_tx_req_only_maint_req): LOG MAINT only transmits MAINT requests

  //*COVERAGE*
  //(cp_tx_req_arb_stall_mid_packet): The arbiter stalls the LOG Maint mid-request
  //(cp_tx_req_arb_stall_btw_packets): The arbiter stalls the LOG Maint between requests
  //(cp_tx_req_arb_stall_first_beat): The arbiter stalls the LOG Maint on the first beat of a request

  // }}} end Arbiter Request Interface - lrq

  endmodule

// {{{ DISCLAIMER OF LIABILITY
// -----------------------------------------------------------------
// (c) Copyright 2011-2013 Xilinx, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
// }}}




//protect end

